library verilog;
use verilog.vl_types.all;
entity altera_avalon_mm_master_bfm is
    generic(
        AV_ADDRESS_W    : integer := 32;
        AV_SYMBOL_W     : integer := 8;
        AV_NUMSYMBOLS   : integer := 4;
        AV_BURSTCOUNT_W : integer := 3;
        AV_READRESPONSE_W: integer := 8;
        AV_WRITERESPONSE_W: integer := 8;
        USE_READ        : integer := 1;
        USE_WRITE       : integer := 1;
        USE_ADDRESS     : integer := 1;
        USE_BYTE_ENABLE : integer := 1;
        USE_BURSTCOUNT  : integer := 1;
        USE_READ_DATA   : integer := 1;
        USE_READ_DATA_VALID: integer := 1;
        USE_WRITE_DATA  : integer := 1;
        USE_BEGIN_TRANSFER: integer := 1;
        USE_BEGIN_BURST_TRANSFER: integer := 1;
        USE_WAIT_REQUEST: integer := 1;
        USE_ARBITERLOCK : integer := 0;
        USE_LOCK        : integer := 0;
        USE_DEBUGACCESS : integer := 0;
        USE_TRANSACTIONID: integer := 0;
        USE_WRITERESPONSE: integer := 0;
        USE_READRESPONSE: integer := 0;
        USE_CLKEN       : integer := 0;
        AV_REGISTERINCOMINGSIGNALS: integer := 0;
        AV_FIX_READ_LATENCY: integer := 0;
        AV_MAX_PENDING_READS: integer := 0;
        AV_MAX_PENDING_WRITES: integer := 0;
        AV_BURST_LINEWRAP: integer := 0;
        AV_BURST_BNDR_ONLY: integer := 0;
        AV_CONSTANT_BURST_BEHAVIOR: integer := 1;
        AV_READ_WAIT_TIME: integer := 0;
        AV_WRITE_WAIT_TIME: integer := 0;
        REGISTER_WAITREQUEST: integer := 0;
        VHDL_ID         : integer := 0
    );
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        avm_clken       : out    vl_logic;
        avm_waitrequest : in     vl_logic;
        avm_write       : out    vl_logic;
        avm_read        : out    vl_logic;
        avm_address     : out    vl_logic_vector;
        avm_byteenable  : out    vl_logic_vector;
        avm_burstcount  : out    vl_logic_vector;
        avm_beginbursttransfer: out    vl_logic;
        avm_begintransfer: out    vl_logic;
        avm_writedata   : out    vl_logic_vector;
        avm_readdata    : in     vl_logic_vector;
        avm_readdatavalid: in     vl_logic;
        avm_arbiterlock : out    vl_logic;
        avm_lock        : out    vl_logic;
        avm_debugaccess : out    vl_logic;
        avm_transactionid: out    vl_logic_vector(7 downto 0);
        avm_readresponse: in     vl_logic_vector;
        avm_readid      : in     vl_logic_vector(7 downto 0);
        avm_writeresponserequest: out    vl_logic;
        avm_writeresponsevalid: in     vl_logic;
        avm_writeresponse: in     vl_logic_vector;
        avm_writeid     : in     vl_logic_vector(7 downto 0);
        avm_response    : in     vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AV_ADDRESS_W : constant is 1;
    attribute mti_svvh_generic_type of AV_SYMBOL_W : constant is 1;
    attribute mti_svvh_generic_type of AV_NUMSYMBOLS : constant is 1;
    attribute mti_svvh_generic_type of AV_BURSTCOUNT_W : constant is 1;
    attribute mti_svvh_generic_type of AV_READRESPONSE_W : constant is 1;
    attribute mti_svvh_generic_type of AV_WRITERESPONSE_W : constant is 1;
    attribute mti_svvh_generic_type of USE_READ : constant is 1;
    attribute mti_svvh_generic_type of USE_WRITE : constant is 1;
    attribute mti_svvh_generic_type of USE_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of USE_BYTE_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of USE_BURSTCOUNT : constant is 1;
    attribute mti_svvh_generic_type of USE_READ_DATA : constant is 1;
    attribute mti_svvh_generic_type of USE_READ_DATA_VALID : constant is 1;
    attribute mti_svvh_generic_type of USE_WRITE_DATA : constant is 1;
    attribute mti_svvh_generic_type of USE_BEGIN_TRANSFER : constant is 1;
    attribute mti_svvh_generic_type of USE_BEGIN_BURST_TRANSFER : constant is 1;
    attribute mti_svvh_generic_type of USE_WAIT_REQUEST : constant is 1;
    attribute mti_svvh_generic_type of USE_ARBITERLOCK : constant is 1;
    attribute mti_svvh_generic_type of USE_LOCK : constant is 1;
    attribute mti_svvh_generic_type of USE_DEBUGACCESS : constant is 1;
    attribute mti_svvh_generic_type of USE_TRANSACTIONID : constant is 1;
    attribute mti_svvh_generic_type of USE_WRITERESPONSE : constant is 1;
    attribute mti_svvh_generic_type of USE_READRESPONSE : constant is 1;
    attribute mti_svvh_generic_type of USE_CLKEN : constant is 1;
    attribute mti_svvh_generic_type of AV_REGISTERINCOMINGSIGNALS : constant is 1;
    attribute mti_svvh_generic_type of AV_FIX_READ_LATENCY : constant is 1;
    attribute mti_svvh_generic_type of AV_MAX_PENDING_READS : constant is 1;
    attribute mti_svvh_generic_type of AV_MAX_PENDING_WRITES : constant is 1;
    attribute mti_svvh_generic_type of AV_BURST_LINEWRAP : constant is 1;
    attribute mti_svvh_generic_type of AV_BURST_BNDR_ONLY : constant is 1;
    attribute mti_svvh_generic_type of AV_CONSTANT_BURST_BEHAVIOR : constant is 1;
    attribute mti_svvh_generic_type of AV_READ_WAIT_TIME : constant is 1;
    attribute mti_svvh_generic_type of AV_WRITE_WAIT_TIME : constant is 1;
    attribute mti_svvh_generic_type of REGISTER_WAITREQUEST : constant is 1;
    attribute mti_svvh_generic_type of VHDL_ID : constant is 1;
end altera_avalon_mm_master_bfm;
