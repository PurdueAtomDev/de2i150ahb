library verilog;
use verilog.vl_types.all;
entity cycloneiv_hssi_tx_digi is
    port(
        txpcs_rst       : in     vl_logic;
        scan_mode       : in     vl_logic;
        txd             : in     vl_logic_vector(43 downto 0);
        pld_tx_clk      : in     vl_logic;
        polinv_tx       : in     vl_logic;
        rev_loop_data   : in     vl_logic_vector(19 downto 0);
        wrenable_tx     : in     vl_logic;
        rddisable_tx    : in     vl_logic;
        phfifourst_tx   : in     vl_logic;
        txdetectrxloopback: in     vl_logic;
        powerdown       : in     vl_logic_vector(1 downto 0);
        revloopback     : in     vl_logic;
        txswing         : in     vl_logic;
        pcs_txdeemph    : in     vl_logic;
        pcs_txmargin    : in     vl_logic_vector(2 downto 0);
        rxpolarity      : in     vl_logic;
        polinv_rx       : in     vl_logic;
        full_tx         : out    vl_logic;
        empty_tx        : out    vl_logic;
        tx_data_ts      : in     vl_logic_vector(7 downto 0);
        tx_ctl_ts       : in     vl_logic;
        refclk_pma      : in     vl_logic;
        txpma_local_clk : in     vl_logic;
        tx_clk_out      : out    vl_logic;
        tx_data_tc      : out    vl_logic_vector(7 downto 0);
        tx_ctl_tc       : out    vl_logic;
        pudr            : out    vl_logic_vector(19 downto 0);
        rd_enable_sync  : out    vl_logic;
        refclk_b        : out    vl_logic;
        txlp20b         : out    vl_logic_vector(19 downto 0);
        tx_pipe_clk     : out    vl_logic;
        encoder_testbus : out    vl_logic_vector(9 downto 0);
        tx_ctrl_testbus : out    vl_logic_vector(9 downto 0);
        tx_pipe_soft_reset: out    vl_logic;
        tx_pipe_electidle: out    vl_logic;
        txdetectrxloopback_int: out    vl_logic;
        powerdown_int   : out    vl_logic_vector(1 downto 0);
        revloopback_int : out    vl_logic;
        phfifo_txswing  : out    vl_logic;
        phfifo_txdeemph : out    vl_logic;
        phfifo_txmargin : out    vl_logic_vector(2 downto 0);
        rxpolarity_int  : out    vl_logic;
        polinv_rx_int   : out    vl_logic;
        rrev_loopbk     : in     vl_logic;
        rev_loopbk      : in     vl_logic;
        eidleinfersel   : in     vl_logic_vector(2 downto 0);
        gray_eidleinfersel: out    vl_logic_vector(2 downto 0);
        rbisten_tx      : in     vl_logic;
        rforce_disp     : in     vl_logic;
        rib_force_disp  : in     vl_logic;
        rforce_echar    : in     vl_logic;
        rforce_kchar    : in     vl_logic;
        rendec_tx       : in     vl_logic;
        rge_xaui_tx     : in     vl_logic;
        rdwidth_tx      : in     vl_logic;
        rtxfifo_dis     : in     vl_logic;
        rcascaded_8b10b_en_tx: in     vl_logic;
        rprbsen_tx      : in     vl_logic;
        rprbs_sel       : in     vl_logic_vector(2 downto 0);
        rbist_sel       : in     vl_logic_vector(1 downto 0);
        rcxpat_chnl_en  : in     vl_logic_vector(1 downto 0);
        renpolinv_tx    : in     vl_logic;
        rphfifopldentx  : in     vl_logic;
        rphfifoursttx   : in     vl_logic;
        rfreerun_tx     : in     vl_logic;
        rtxwrclksel     : in     vl_logic;
        rtxrdclksel     : in     vl_logic;
        renbitrev_tx    : in     vl_logic;
        rensymswap_tx   : in     vl_logic;
        r8b10b_enc_ibm_en: in     vl_logic;
        rtxfifo_lowlatency_en: in     vl_logic;
        rpmadwidth_tx   : in     vl_logic;
        rpma_doublewidth_tx: in     vl_logic;
        rtx_pipe_enable : in     vl_logic;
        rindv_tx        : in     vl_logic;
        rendec_data_sel_tx: in     vl_logic;
        rtxpcsbypass_en : in     vl_logic;
        rtxpcsclkpwdn   : in     vl_logic;
        rauto_speed_ena : in     vl_logic;
        rfreq_sel       : in     vl_logic;
        gen2ngen1       : in     vl_logic;
        gen2ngen1_bundle: in     vl_logic;
        rcid_pattern_tx : in     vl_logic;
        rcid_len_tx     : in     vl_logic_vector(7 downto 0);
        tx_div2_sync_in_centrl: in     vl_logic;
        tx_div2_sync_in_quad_up: in     vl_logic;
        tx_div2_sync_in_quad_down: in     vl_logic;
        wr_enable_in_centrl: in     vl_logic;
        wr_enable_in_quad_up: in     vl_logic;
        wr_enable_in_quad_down: in     vl_logic;
        rd_enable_in_centrl: in     vl_logic;
        rd_enable_in_quad_up: in     vl_logic;
        rd_enable_in_quad_down: in     vl_logic;
        fifo_select_in_centrl: in     vl_logic;
        fifo_select_in_quad_up: in     vl_logic;
        fifo_select_in_quad_down: in     vl_logic;
        dis_pc_byte     : in     vl_logic;
        reset_pc_ptrs   : in     vl_logic;
        reset_pc_ptrs_in_centrl: in     vl_logic;
        reset_pc_ptrs_in_quad_up: in     vl_logic;
        reset_pc_ptrs_in_quad_down: in     vl_logic;
        tx_div2_sync_in_pipe_quad_up: in     vl_logic;
        tx_div2_sync_in_pipe_quad_down: in     vl_logic;
        wr_enable_in_pipe_quad_up: in     vl_logic;
        wr_enable_in_pipe_quad_down: in     vl_logic;
        rd_enable_in_pipe_quad_up: in     vl_logic;
        rd_enable_in_pipe_quad_down: in     vl_logic;
        fifo_select_in_pipe_quad_up: in     vl_logic;
        fifo_select_in_pipe_quad_down: in     vl_logic;
        rmaster_tx      : in     vl_logic;
        rmaster_up_tx   : in     vl_logic;
        rself_sw_en_tx  : in     vl_logic;
        rpipeline_bypass_tx: in     vl_logic;
        rphfifo_regmode_tx: in     vl_logic;
        rtxbitslip_en   : in     vl_logic;
        tx_div2_sync_out_pipe_up: out    vl_logic;
        fifo_select_out_pipe_up: out    vl_logic;
        wr_enable_out_pipe_up: out    vl_logic;
        rd_enable_out_pipe_up: out    vl_logic;
        tx_div2_sync_out_pipe_down: out    vl_logic;
        fifo_select_out_pipe_down: out    vl_logic;
        wr_enable_out_pipe_down: out    vl_logic;
        rd_enable_out_pipe_down: out    vl_logic;
        prbs_cid_en     : in     vl_logic;
        tx_boundary_sel : in     vl_logic_vector(4 downto 0)
    );
end cycloneiv_hssi_tx_digi;
