// ahb_master_slave_with_qsys_bfm.v

// Generated using ACDS version 14.0 200 at 2015.08.10.14:24:38

`timescale 1 ps / 1 ps
module ahb_master_slave_with_qsys_bfm (
		input  wire        clk_clk,                                       //                              clk.clk
		input  wire        reset_reset_n,                                 //                            reset.reset_n
		input  wire        ahb_master_slave_2_0_conduit_end_add_data_sel, // ahb_master_slave_2_0_conduit_end.add_data_sel
		output wire [31:0] ahb_master_slave_2_0_conduit_end_display_data, //                                 .display_data
		input  wire [15:0] ahb_master_slave_2_0_conduit_end_rdwr_address  //                                 .rdwr_address
	);

	wire         avalon2ahb_bridge_0_ahb_master_hwrite;                            // avalon2ahb_bridge_0:HWRITE -> ahb_master_slave_2_0:slave_HWRITE
	wire  [31:0] avalon2ahb_bridge_0_ahb_master_hwdata;                            // avalon2ahb_bridge_0:HWDATA -> ahb_master_slave_2_0:slave_HWDATA
	wire   [3:0] avalon2ahb_bridge_0_ahb_master_hprot;                             // avalon2ahb_bridge_0:HPROT -> ahb_master_slave_2_0:slave_HPROT
	wire         avalon2ahb_bridge_0_ahb_master_hreadyin;                          // avalon2ahb_bridge_0:HREADYIN -> ahb_master_slave_2_0:slave_HREADY
	wire   [2:0] avalon2ahb_bridge_0_ahb_master_hsize;                             // avalon2ahb_bridge_0:HSIZE -> ahb_master_slave_2_0:slave_HSIZE
	wire  [31:0] avalon2ahb_bridge_0_ahb_master_hrdata;                            // ahb_master_slave_2_0:slave_HRDATA -> avalon2ahb_bridge_0:HRDATA
	wire         avalon2ahb_bridge_0_ahb_master_hsel;                              // avalon2ahb_bridge_0:HSEL -> ahb_master_slave_2_0:slave_HSEL
	wire   [1:0] avalon2ahb_bridge_0_ahb_master_htrans;                            // avalon2ahb_bridge_0:HTRANS -> ahb_master_slave_2_0:slave_HTRANS
	wire   [1:0] avalon2ahb_bridge_0_ahb_master_hresp;                             // ahb_master_slave_2_0:slave_HRESP -> avalon2ahb_bridge_0:HRESP
	wire  [31:0] avalon2ahb_bridge_0_ahb_master_haddr;                             // avalon2ahb_bridge_0:HADDR -> ahb_master_slave_2_0:slave_HADDR
	wire         avalon2ahb_bridge_0_ahb_master_hready;                            // ahb_master_slave_2_0:slave_HREADYOUT -> avalon2ahb_bridge_0:HREADY
	wire   [2:0] avalon2ahb_bridge_0_ahb_master_hburst;                            // avalon2ahb_bridge_0:HBURST -> ahb_master_slave_2_0:slave_HBURST
	wire         ahb_master_slave_2_0_ahb_master_hwrite;                           // ahb_master_slave_2_0:master_HWRITE -> ahb2avalon_burst_bridge_0:HWRITE
	wire  [31:0] ahb_master_slave_2_0_ahb_master_hwdata;                           // ahb_master_slave_2_0:master_HWDATA -> ahb2avalon_burst_bridge_0:HWDATA
	wire   [3:0] ahb_master_slave_2_0_ahb_master_hprot;                            // ahb_master_slave_2_0:master_HPROT -> ahb2avalon_burst_bridge_0:HPROT
	wire         ahb_master_slave_2_0_ahb_master_hreadyin;                         // ahb_master_slave_2_0:master_HREADYIN -> ahb2avalon_burst_bridge_0:HREADY
	wire   [2:0] ahb_master_slave_2_0_ahb_master_hsize;                            // ahb_master_slave_2_0:master_HSIZE -> ahb2avalon_burst_bridge_0:HSIZE
	wire  [31:0] ahb_master_slave_2_0_ahb_master_hrdata;                           // ahb2avalon_burst_bridge_0:HRDATA -> ahb_master_slave_2_0:master_HRDATA
	wire         ahb_master_slave_2_0_ahb_master_hsel;                             // ahb_master_slave_2_0:master_HSEL -> ahb2avalon_burst_bridge_0:HSEL
	wire   [1:0] ahb_master_slave_2_0_ahb_master_htrans;                           // ahb_master_slave_2_0:master_HTRANS -> ahb2avalon_burst_bridge_0:HTRANS
	wire   [1:0] ahb_master_slave_2_0_ahb_master_hresp;                            // ahb2avalon_burst_bridge_0:HRESP -> ahb_master_slave_2_0:master_HRESP
	wire         ahb_master_slave_2_0_ahb_master_hready;                           // ahb2avalon_burst_bridge_0:HREADYOUT -> ahb_master_slave_2_0:master_HREADY
	wire  [31:0] ahb_master_slave_2_0_ahb_master_haddr;                            // ahb_master_slave_2_0:master_HADDR -> ahb2avalon_burst_bridge_0:HADDR
	wire   [2:0] ahb_master_slave_2_0_ahb_master_hburst;                           // ahb_master_slave_2_0:master_HBURST -> ahb2avalon_burst_bridge_0:HBURST
	wire         mm_master_bfm_0_m0_waitrequest;                                   // mm_interconnect_0:mm_master_bfm_0_m0_waitrequest -> mm_master_bfm_0:avm_waitrequest
	wire   [2:0] mm_master_bfm_0_m0_burstcount;                                    // mm_master_bfm_0:avm_burstcount -> mm_interconnect_0:mm_master_bfm_0_m0_burstcount
	wire  [31:0] mm_master_bfm_0_m0_writedata;                                     // mm_master_bfm_0:avm_writedata -> mm_interconnect_0:mm_master_bfm_0_m0_writedata
	wire  [31:0] mm_master_bfm_0_m0_address;                                       // mm_master_bfm_0:avm_address -> mm_interconnect_0:mm_master_bfm_0_m0_address
	wire         mm_master_bfm_0_m0_write;                                         // mm_master_bfm_0:avm_write -> mm_interconnect_0:mm_master_bfm_0_m0_write
	wire         mm_master_bfm_0_m0_read;                                          // mm_master_bfm_0:avm_read -> mm_interconnect_0:mm_master_bfm_0_m0_read
	wire  [31:0] mm_master_bfm_0_m0_readdata;                                      // mm_interconnect_0:mm_master_bfm_0_m0_readdata -> mm_master_bfm_0:avm_readdata
	wire         mm_master_bfm_0_m0_readdatavalid;                                 // mm_interconnect_0:mm_master_bfm_0_m0_readdatavalid -> mm_master_bfm_0:avm_readdatavalid
	wire   [3:0] mm_master_bfm_0_m0_byteenable;                                    // mm_master_bfm_0:avm_byteenable -> mm_interconnect_0:mm_master_bfm_0_m0_byteenable
	wire         mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_waitrequest;   // avalon2ahb_bridge_0:waitrequest -> mm_interconnect_0:avalon2ahb_bridge_0_avalon_slave_waitrequest
	wire  [31:0] mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_writedata;     // mm_interconnect_0:avalon2ahb_bridge_0_avalon_slave_writedata -> avalon2ahb_bridge_0:writedata
	wire   [4:0] mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_address;       // mm_interconnect_0:avalon2ahb_bridge_0_avalon_slave_address -> avalon2ahb_bridge_0:address
	wire         mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_write;         // mm_interconnect_0:avalon2ahb_bridge_0_avalon_slave_write -> avalon2ahb_bridge_0:write
	wire         mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_read;          // mm_interconnect_0:avalon2ahb_bridge_0_avalon_slave_read -> avalon2ahb_bridge_0:read
	wire  [31:0] mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_readdata;      // avalon2ahb_bridge_0:readdata -> mm_interconnect_0:avalon2ahb_bridge_0_avalon_slave_readdata
	wire         mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_readdatavalid; // avalon2ahb_bridge_0:readdatavalid -> mm_interconnect_0:avalon2ahb_bridge_0_avalon_slave_readdatavalid
	wire   [3:0] ahb2avalon_burst_bridge_0_avalon_master_burstcount;               // ahb2avalon_burst_bridge_0:burstcount -> mm_interconnect_3:ahb2avalon_burst_bridge_0_avalon_master_burstcount
	wire         ahb2avalon_burst_bridge_0_avalon_master_waitrequest;              // mm_interconnect_3:ahb2avalon_burst_bridge_0_avalon_master_waitrequest -> ahb2avalon_burst_bridge_0:waitrequest
	wire  [31:0] ahb2avalon_burst_bridge_0_avalon_master_writedata;                // ahb2avalon_burst_bridge_0:writedata -> mm_interconnect_3:ahb2avalon_burst_bridge_0_avalon_master_writedata
	wire  [31:0] ahb2avalon_burst_bridge_0_avalon_master_address;                  // ahb2avalon_burst_bridge_0:address -> mm_interconnect_3:ahb2avalon_burst_bridge_0_avalon_master_address
	wire         ahb2avalon_burst_bridge_0_avalon_master_write;                    // ahb2avalon_burst_bridge_0:write -> mm_interconnect_3:ahb2avalon_burst_bridge_0_avalon_master_write
	wire         ahb2avalon_burst_bridge_0_avalon_master_read;                     // ahb2avalon_burst_bridge_0:read -> mm_interconnect_3:ahb2avalon_burst_bridge_0_avalon_master_read
	wire  [31:0] ahb2avalon_burst_bridge_0_avalon_master_readdata;                 // mm_interconnect_3:ahb2avalon_burst_bridge_0_avalon_master_readdata -> ahb2avalon_burst_bridge_0:readdata
	wire         ahb2avalon_burst_bridge_0_avalon_master_readdatavalid;            // mm_interconnect_3:ahb2avalon_burst_bridge_0_avalon_master_readdatavalid -> ahb2avalon_burst_bridge_0:readdatavalid
	wire   [3:0] ahb2avalon_burst_bridge_0_avalon_master_byteenable;               // ahb2avalon_burst_bridge_0:byteenable -> mm_interconnect_3:ahb2avalon_burst_bridge_0_avalon_master_byteenable
	wire         mm_interconnect_3_mm_slave_bfm_0_s0_waitrequest;                  // mm_slave_bfm_0:avs_waitrequest -> mm_interconnect_3:mm_slave_bfm_0_s0_waitrequest
	wire  [31:0] mm_interconnect_3_mm_slave_bfm_0_s0_writedata;                    // mm_interconnect_3:mm_slave_bfm_0_s0_writedata -> mm_slave_bfm_0:avs_writedata
	wire   [4:0] mm_interconnect_3_mm_slave_bfm_0_s0_address;                      // mm_interconnect_3:mm_slave_bfm_0_s0_address -> mm_slave_bfm_0:avs_address
	wire         mm_interconnect_3_mm_slave_bfm_0_s0_write;                        // mm_interconnect_3:mm_slave_bfm_0_s0_write -> mm_slave_bfm_0:avs_write
	wire         mm_interconnect_3_mm_slave_bfm_0_s0_read;                         // mm_interconnect_3:mm_slave_bfm_0_s0_read -> mm_slave_bfm_0:avs_read
	wire  [31:0] mm_interconnect_3_mm_slave_bfm_0_s0_readdata;                     // mm_slave_bfm_0:avs_readdata -> mm_interconnect_3:mm_slave_bfm_0_s0_readdata
	wire         mm_interconnect_3_mm_slave_bfm_0_s0_readdatavalid;                // mm_slave_bfm_0:avs_readdatavalid -> mm_interconnect_3:mm_slave_bfm_0_s0_readdatavalid
	wire   [3:0] mm_interconnect_3_mm_slave_bfm_0_s0_byteenable;                   // mm_interconnect_3:mm_slave_bfm_0_s0_byteenable -> mm_slave_bfm_0:avs_byteenable
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [ahb2avalon_burst_bridge_0:reset_n, ahb_master_slave_2_0:HRESETn, avalon2ahb_bridge_0:reset_n, mm_interconnect_0:mm_master_bfm_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_3:ahb2avalon_burst_bridge_0_reset_reset_bridge_in_reset_reset, mm_master_bfm_0:reset, mm_slave_bfm_0:reset]

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (32),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) mm_master_bfm_0 (
		.clk                      (clk_clk),                          //       clk.clk
		.reset                    (rst_controller_reset_out_reset),   // clk_reset.reset
		.avm_address              (mm_master_bfm_0_m0_address),       //        m0.address
		.avm_burstcount           (mm_master_bfm_0_m0_burstcount),    //          .burstcount
		.avm_readdata             (mm_master_bfm_0_m0_readdata),      //          .readdata
		.avm_writedata            (mm_master_bfm_0_m0_writedata),     //          .writedata
		.avm_waitrequest          (mm_master_bfm_0_m0_waitrequest),   //          .waitrequest
		.avm_write                (mm_master_bfm_0_m0_write),         //          .write
		.avm_read                 (mm_master_bfm_0_m0_read),          //          .read
		.avm_byteenable           (mm_master_bfm_0_m0_byteenable),    //          .byteenable
		.avm_readdatavalid        (mm_master_bfm_0_m0_readdatavalid), //          .readdatavalid
		.avm_begintransfer        (),                                 // (terminated)
		.avm_beginbursttransfer   (),                                 // (terminated)
		.avm_arbiterlock          (),                                 // (terminated)
		.avm_lock                 (),                                 // (terminated)
		.avm_debugaccess          (),                                 // (terminated)
		.avm_transactionid        (),                                 // (terminated)
		.avm_readid               (8'b00000000),                      // (terminated)
		.avm_writeid              (8'b00000000),                      // (terminated)
		.avm_clken                (),                                 // (terminated)
		.avm_response             (2'b00),                            // (terminated)
		.avm_writeresponserequest (),                                 // (terminated)
		.avm_writeresponsevalid   (1'b0),                             // (terminated)
		.avm_readresponse         (8'b00000000),                      // (terminated)
		.avm_writeresponse        (8'b00000000)                       // (terminated)
	);

	altera_avalon_mm_slave_bfm #(
		.AV_ADDRESS_W               (5),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (4),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (32),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) mm_slave_bfm_0 (
		.clk                      (clk_clk),                                           //       clk.clk
		.reset                    (rst_controller_reset_out_reset),                    // clk_reset.reset
		.avs_writedata            (mm_interconnect_3_mm_slave_bfm_0_s0_writedata),     //        s0.writedata
		.avs_readdata             (mm_interconnect_3_mm_slave_bfm_0_s0_readdata),      //          .readdata
		.avs_address              (mm_interconnect_3_mm_slave_bfm_0_s0_address),       //          .address
		.avs_waitrequest          (mm_interconnect_3_mm_slave_bfm_0_s0_waitrequest),   //          .waitrequest
		.avs_write                (mm_interconnect_3_mm_slave_bfm_0_s0_write),         //          .write
		.avs_read                 (mm_interconnect_3_mm_slave_bfm_0_s0_read),          //          .read
		.avs_byteenable           (mm_interconnect_3_mm_slave_bfm_0_s0_byteenable),    //          .byteenable
		.avs_readdatavalid        (mm_interconnect_3_mm_slave_bfm_0_s0_readdatavalid), //          .readdatavalid
		.avs_begintransfer        (1'b0),                                              // (terminated)
		.avs_beginbursttransfer   (1'b0),                                              // (terminated)
		.avs_burstcount           (4'b0001),                                           // (terminated)
		.avs_arbiterlock          (1'b0),                                              // (terminated)
		.avs_lock                 (1'b0),                                              // (terminated)
		.avs_debugaccess          (1'b0),                                              // (terminated)
		.avs_transactionid        (8'b00000000),                                       // (terminated)
		.avs_readid               (),                                                  // (terminated)
		.avs_writeid              (),                                                  // (terminated)
		.avs_clken                (1'b1),                                              // (terminated)
		.avs_response             (),                                                  // (terminated)
		.avs_writeresponserequest (1'b0),                                              // (terminated)
		.avs_writeresponsevalid   (),                                                  // (terminated)
		.avs_readresponse         (),                                                  // (terminated)
		.avs_writeresponse        ()                                                   // (terminated)
	);

	top_level ahb_master_slave_2_0 (
		.add_data_sel    (ahb_master_slave_2_0_conduit_end_add_data_sel), // conduit_end.add_data_sel
		.display_data    (ahb_master_slave_2_0_conduit_end_display_data), //            .display_data
		.rdwr_address    (ahb_master_slave_2_0_conduit_end_rdwr_address), //            .rdwr_address
		.HRESETn         (~rst_controller_reset_out_reset),               //  reset_sink.reset_n
		.HCLK            (clk_clk),                                       //  clock_sink.clk
		.slave_HADDR     (avalon2ahb_bridge_0_ahb_master_haddr),          //   ahb_slave.haddr
		.slave_HBURST    (avalon2ahb_bridge_0_ahb_master_hburst),         //            .hburst
		.slave_HPROT     (avalon2ahb_bridge_0_ahb_master_hprot),          //            .hprot
		.slave_HSIZE     (avalon2ahb_bridge_0_ahb_master_hsize),          //            .hsize
		.slave_HTRANS    (avalon2ahb_bridge_0_ahb_master_htrans),         //            .htrans
		.slave_HWDATA    (avalon2ahb_bridge_0_ahb_master_hwdata),         //            .hwdata
		.slave_HWRITE    (avalon2ahb_bridge_0_ahb_master_hwrite),         //            .hwrite
		.slave_HRDATA    (avalon2ahb_bridge_0_ahb_master_hrdata),         //            .hrdata
		.slave_HREADYOUT (avalon2ahb_bridge_0_ahb_master_hready),         //            .hready
		.slave_HRESP     (avalon2ahb_bridge_0_ahb_master_hresp),          //            .hresp
		.slave_HSEL      (avalon2ahb_bridge_0_ahb_master_hsel),           //            .hsel
		.slave_HREADY    (avalon2ahb_bridge_0_ahb_master_hreadyin),       //            .hreadyin
		.master_HADDR    (ahb_master_slave_2_0_ahb_master_haddr),         //  ahb_master.haddr
		.master_HBURST   (ahb_master_slave_2_0_ahb_master_hburst),        //            .hburst
		.master_HPROT    (ahb_master_slave_2_0_ahb_master_hprot),         //            .hprot
		.master_HSIZE    (ahb_master_slave_2_0_ahb_master_hsize),         //            .hsize
		.master_HTRANS   (ahb_master_slave_2_0_ahb_master_htrans),        //            .htrans
		.master_HWDATA   (ahb_master_slave_2_0_ahb_master_hwdata),        //            .hwdata
		.master_HWRITE   (ahb_master_slave_2_0_ahb_master_hwrite),        //            .hwrite
		.master_HRDATA   (ahb_master_slave_2_0_ahb_master_hrdata),        //            .hrdata
		.master_HREADY   (ahb_master_slave_2_0_ahb_master_hready),        //            .hready
		.master_HRESP    (ahb_master_slave_2_0_ahb_master_hresp),         //            .hresp
		.master_HREADYIN (ahb_master_slave_2_0_ahb_master_hreadyin),      //            .hreadyin
		.master_HSEL     (ahb_master_slave_2_0_ahb_master_hsel)           //            .hsel
	);

	avalon_ahb_bridge #(
		.AVALON_ADDRESSWIDTH (5),
		.ADDRESSWIDTH        (32),
		.DATAWIDTH           (32)
	) avalon2ahb_bridge_0 (
		.clk           (clk_clk),                                                          //        clock.clk
		.reset_n       (~rst_controller_reset_out_reset),                                  //        reset.reset_n
		.read          (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_read),          // avalon_slave.read
		.address       (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_address),       //             .address
		.write         (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_write),         //             .write
		.writedata     (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_writedata),     //             .writedata
		.waitrequest   (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_waitrequest),   //             .waitrequest
		.readdatavalid (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_readdatavalid), //             .readdatavalid
		.readdata      (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_readdata),      //             .readdata
		.HRDATA        (avalon2ahb_bridge_0_ahb_master_hrdata),                            //   ahb_master.hrdata
		.HREADY        (avalon2ahb_bridge_0_ahb_master_hready),                            //             .hready
		.HRESP         (avalon2ahb_bridge_0_ahb_master_hresp),                             //             .hresp
		.HBURST        (avalon2ahb_bridge_0_ahb_master_hburst),                            //             .hburst
		.HSIZE         (avalon2ahb_bridge_0_ahb_master_hsize),                             //             .hsize
		.HTRANS        (avalon2ahb_bridge_0_ahb_master_htrans),                            //             .htrans
		.HSEL          (avalon2ahb_bridge_0_ahb_master_hsel),                              //             .hsel
		.HPROT         (avalon2ahb_bridge_0_ahb_master_hprot),                             //             .hprot
		.HADDR         (avalon2ahb_bridge_0_ahb_master_haddr),                             //             .haddr
		.HWDATA        (avalon2ahb_bridge_0_ahb_master_hwdata),                            //             .hwdata
		.HWRITE        (avalon2ahb_bridge_0_ahb_master_hwrite),                            //             .hwrite
		.HREADYIN      (avalon2ahb_bridge_0_ahb_master_hreadyin)                           //             .hreadyin
	);

	ahb_avalon_bridge_with_burst #(
		.ADDRESSWIDTH  (32),
		.DATAWIDTH     (32),
		.FIFODEPTH     (32),
		.FIFODEPTH_LOG (5),
		.MAXBURSTCOUNT (8)
	) ahb2avalon_burst_bridge_0 (
		.clk           (clk_clk),                                               //         clock.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.address       (ahb2avalon_burst_bridge_0_avalon_master_address),       // avalon_master.address
		.write         (ahb2avalon_burst_bridge_0_avalon_master_write),         //              .write
		.read          (ahb2avalon_burst_bridge_0_avalon_master_read),          //              .read
		.byteenable    (ahb2avalon_burst_bridge_0_avalon_master_byteenable),    //              .byteenable
		.writedata     (ahb2avalon_burst_bridge_0_avalon_master_writedata),     //              .writedata
		.waitrequest   (ahb2avalon_burst_bridge_0_avalon_master_waitrequest),   //              .waitrequest
		.readdatavalid (ahb2avalon_burst_bridge_0_avalon_master_readdatavalid), //              .readdatavalid
		.readdata      (ahb2avalon_burst_bridge_0_avalon_master_readdata),      //              .readdata
		.burstcount    (ahb2avalon_burst_bridge_0_avalon_master_burstcount),    //              .burstcount
		.HRDATA        (ahb_master_slave_2_0_ahb_master_hrdata),                //     ahb_slave.hrdata
		.HREADY        (ahb_master_slave_2_0_ahb_master_hreadyin),              //              .hreadyin
		.HRESP         (ahb_master_slave_2_0_ahb_master_hresp),                 //              .hresp
		.HBURST        (ahb_master_slave_2_0_ahb_master_hburst),                //              .hburst
		.HSIZE         (ahb_master_slave_2_0_ahb_master_hsize),                 //              .hsize
		.HTRANS        (ahb_master_slave_2_0_ahb_master_htrans),                //              .htrans
		.HPROT         (ahb_master_slave_2_0_ahb_master_hprot),                 //              .hprot
		.HADDR         (ahb_master_slave_2_0_ahb_master_haddr),                 //              .haddr
		.HWDATA        (ahb_master_slave_2_0_ahb_master_hwdata),                //              .hwdata
		.HWRITE        (ahb_master_slave_2_0_ahb_master_hwrite),                //              .hwrite
		.HREADYOUT     (ahb_master_slave_2_0_ahb_master_hready),                //              .hready
		.HSEL          (ahb_master_slave_2_0_ahb_master_hsel)                   //              .hsel
	);

	ahb_master_slave_with_qsys_bfm_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                         (clk_clk),                                                          //                                       clk_0_clk.clk
		.mm_master_bfm_0_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                   // mm_master_bfm_0_clk_reset_reset_bridge_in_reset.reset
		.mm_master_bfm_0_m0_address                            (mm_master_bfm_0_m0_address),                                       //                              mm_master_bfm_0_m0.address
		.mm_master_bfm_0_m0_waitrequest                        (mm_master_bfm_0_m0_waitrequest),                                   //                                                .waitrequest
		.mm_master_bfm_0_m0_burstcount                         (mm_master_bfm_0_m0_burstcount),                                    //                                                .burstcount
		.mm_master_bfm_0_m0_byteenable                         (mm_master_bfm_0_m0_byteenable),                                    //                                                .byteenable
		.mm_master_bfm_0_m0_read                               (mm_master_bfm_0_m0_read),                                          //                                                .read
		.mm_master_bfm_0_m0_readdata                           (mm_master_bfm_0_m0_readdata),                                      //                                                .readdata
		.mm_master_bfm_0_m0_readdatavalid                      (mm_master_bfm_0_m0_readdatavalid),                                 //                                                .readdatavalid
		.mm_master_bfm_0_m0_write                              (mm_master_bfm_0_m0_write),                                         //                                                .write
		.mm_master_bfm_0_m0_writedata                          (mm_master_bfm_0_m0_writedata),                                     //                                                .writedata
		.avalon2ahb_bridge_0_avalon_slave_address              (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_address),       //                avalon2ahb_bridge_0_avalon_slave.address
		.avalon2ahb_bridge_0_avalon_slave_write                (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_write),         //                                                .write
		.avalon2ahb_bridge_0_avalon_slave_read                 (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_read),          //                                                .read
		.avalon2ahb_bridge_0_avalon_slave_readdata             (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_readdata),      //                                                .readdata
		.avalon2ahb_bridge_0_avalon_slave_writedata            (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_writedata),     //                                                .writedata
		.avalon2ahb_bridge_0_avalon_slave_readdatavalid        (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_readdatavalid), //                                                .readdatavalid
		.avalon2ahb_bridge_0_avalon_slave_waitrequest          (mm_interconnect_0_avalon2ahb_bridge_0_avalon_slave_waitrequest)    //                                                .waitrequest
	);

	ahb_master_slave_with_qsys_bfm_mm_interconnect_3 mm_interconnect_3 (
		.clk_0_clk_clk                                               (clk_clk),                                               //                                             clk_0_clk.clk
		.ahb2avalon_burst_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // ahb2avalon_burst_bridge_0_reset_reset_bridge_in_reset.reset
		.ahb2avalon_burst_bridge_0_avalon_master_address             (ahb2avalon_burst_bridge_0_avalon_master_address),       //               ahb2avalon_burst_bridge_0_avalon_master.address
		.ahb2avalon_burst_bridge_0_avalon_master_waitrequest         (ahb2avalon_burst_bridge_0_avalon_master_waitrequest),   //                                                      .waitrequest
		.ahb2avalon_burst_bridge_0_avalon_master_burstcount          (ahb2avalon_burst_bridge_0_avalon_master_burstcount),    //                                                      .burstcount
		.ahb2avalon_burst_bridge_0_avalon_master_byteenable          (ahb2avalon_burst_bridge_0_avalon_master_byteenable),    //                                                      .byteenable
		.ahb2avalon_burst_bridge_0_avalon_master_read                (ahb2avalon_burst_bridge_0_avalon_master_read),          //                                                      .read
		.ahb2avalon_burst_bridge_0_avalon_master_readdata            (ahb2avalon_burst_bridge_0_avalon_master_readdata),      //                                                      .readdata
		.ahb2avalon_burst_bridge_0_avalon_master_readdatavalid       (ahb2avalon_burst_bridge_0_avalon_master_readdatavalid), //                                                      .readdatavalid
		.ahb2avalon_burst_bridge_0_avalon_master_write               (ahb2avalon_burst_bridge_0_avalon_master_write),         //                                                      .write
		.ahb2avalon_burst_bridge_0_avalon_master_writedata           (ahb2avalon_burst_bridge_0_avalon_master_writedata),     //                                                      .writedata
		.mm_slave_bfm_0_s0_address                                   (mm_interconnect_3_mm_slave_bfm_0_s0_address),           //                                     mm_slave_bfm_0_s0.address
		.mm_slave_bfm_0_s0_write                                     (mm_interconnect_3_mm_slave_bfm_0_s0_write),             //                                                      .write
		.mm_slave_bfm_0_s0_read                                      (mm_interconnect_3_mm_slave_bfm_0_s0_read),              //                                                      .read
		.mm_slave_bfm_0_s0_readdata                                  (mm_interconnect_3_mm_slave_bfm_0_s0_readdata),          //                                                      .readdata
		.mm_slave_bfm_0_s0_writedata                                 (mm_interconnect_3_mm_slave_bfm_0_s0_writedata),         //                                                      .writedata
		.mm_slave_bfm_0_s0_byteenable                                (mm_interconnect_3_mm_slave_bfm_0_s0_byteenable),        //                                                      .byteenable
		.mm_slave_bfm_0_s0_readdatavalid                             (mm_interconnect_3_mm_slave_bfm_0_s0_readdatavalid),     //                                                      .readdatavalid
		.mm_slave_bfm_0_s0_waitrequest                               (mm_interconnect_3_mm_slave_bfm_0_s0_waitrequest)        //                                                      .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
