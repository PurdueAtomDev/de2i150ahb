library verilog;
use verilog.vl_types.all;
entity cycloneiv_hssi_cmu is
    generic(
        lpm_type        : string  := "cycloneiv_hssi_cmu";
        auto_spd_deassert_ph_fifo_rst_count: integer := 0;
        auto_spd_phystatus_notify_count: integer := 0;
        coreclk_out_gated_by_quad_reset: string  := "false";
        in_xaui_mode    : string  := "false";
        pipe_auto_speed_nego_enable: string  := "false";
        rx_xaui_sm_backward_compatible_enable: string  := "false";
        rx0_channel_bonding: string  := "none";
        rx0_clk1_mux_select: string  := "recovered clock";
        rx0_clk2_mux_select: string  := "recovered clock";
        rx0_clk_pd_enable: string  := "false";
        rx0_ph_fifo_reg_mode: string  := "false";
        rx0_ph_fifo_reset_enable: string  := "false";
        rx0_ph_fifo_user_ctrl_enable: string  := "false";
        rx0_rd_clk_mux_select: string  := "int clock";
        rx0_recovered_clk_mux_select: string  := "recovered clock";
        rx0_reset_clock_output_during_digital_reset: string  := "false";
        rx0_use_double_data_mode: string  := "false";
        select_refclk_dig: string  := "false";
        tx_xaui_sm_backward_compatible_enable: string  := "false";
        tx0_channel_bonding: string  := "none";
        tx0_clk_pd_enable: string  := "false";
        tx0_ph_fifo_reset_enable: string  := "false";
        tx0_ph_fifo_user_ctrl_enable: string  := "false";
        tx0_rd_clk_mux_select: string  := "local";
        tx0_reset_clock_output_during_digital_reset: string  := "false";
        tx0_use_double_data_mode: string  := "false";
        tx0_wr_clk_mux_select: string  := "int_clk";
        use_coreclk_out_post_divider: string  := "false";
        use_deskew_fifo : string  := "false";
        dprio_config_mode: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_logical_to_physical_mapping: integer := -1;
        tx_logical_to_physical_mapping: integer := -1;
        pll_logical_to_physical_mapping: integer := -1;
        portaddr        : integer := 1;
        devaddr         : integer := 1;
        rx0_logical_to_physical_mapping: integer := 0;
        rx1_logical_to_physical_mapping: integer := 1;
        rx2_logical_to_physical_mapping: integer := 2;
        rx3_logical_to_physical_mapping: integer := 3;
        tx0_logical_to_physical_mapping: integer := 0;
        tx1_logical_to_physical_mapping: integer := 1;
        tx2_logical_to_physical_mapping: integer := 2;
        tx3_logical_to_physical_mapping: integer := 3
    );
    port(
        adet            : in     vl_logic_vector(3 downto 0);
        dpclk           : in     vl_logic;
        dpriodisable    : in     vl_logic;
        dprioin         : in     vl_logic;
        dprioload       : in     vl_logic;
        fixedclk        : in     vl_logic_vector(3 downto 0);
        nonuserfromcal  : in     vl_logic;
        pmacramtest     : in     vl_logic;
        quadreset       : in     vl_logic;
        rdalign         : in     vl_logic_vector(3 downto 0);
        recovclk        : in     vl_logic;
        rdenablesync    : in     vl_logic;
        refclkdig       : in     vl_logic;
        rxrunningdisp   : in     vl_logic_vector(3 downto 0);
        rxanalogreset   : in     vl_logic_vector(3 downto 0);
        rxcoreclk       : in     vl_logic;
        rxctrl          : in     vl_logic_vector(3 downto 0);
        rxdatain        : in     vl_logic_vector(31 downto 0);
        rxdatavalid     : in     vl_logic_vector(3 downto 0);
        rxdigitalreset  : in     vl_logic_vector(3 downto 0);
        rxphfifordenable: in     vl_logic;
        rxphfiforeset   : in     vl_logic;
        rxphfifowrdisable: in     vl_logic;
        rxpowerdown     : in     vl_logic_vector(3 downto 0);
        scanclk         : in     vl_logic;
        scanmode        : in     vl_logic;
        scanshift       : in     vl_logic;
        syncstatus      : in     vl_logic_vector(3 downto 0);
        testin          : in     vl_logic_vector(1999 downto 0);
        txclk           : in     vl_logic;
        txcoreclk       : in     vl_logic;
        txctrl          : in     vl_logic_vector(3 downto 0);
        txdatain        : in     vl_logic_vector(31 downto 0);
        txdigitalreset  : in     vl_logic_vector(3 downto 0);
        txphfiforddisable: in     vl_logic;
        txphfiforeset   : in     vl_logic;
        txphfifowrenable: in     vl_logic;
        rxpmadprioin    : in     vl_logic_vector(1199 downto 0);
        rxpcsdprioin    : in     vl_logic_vector(1599 downto 0);
        txpmadprioin    : in     vl_logic_vector(1199 downto 0);
        txpcsdprioin    : in     vl_logic_vector(599 downto 0);
        alignstatus     : out    vl_logic;
        coreclkout      : out    vl_logic;
        digitaltestout  : out    vl_logic_vector(9 downto 0);
        dpriodisableout : out    vl_logic;
        dpriooe         : out    vl_logic;
        dprioout        : out    vl_logic;
        enabledeskew    : out    vl_logic;
        fiforesetrd     : out    vl_logic;
        quadresetout    : out    vl_logic;
        refclkout       : out    vl_logic;
        rxanalogresetout: out    vl_logic_vector(3 downto 0);
        rxcrupowerdown  : out    vl_logic_vector(3 downto 0);
        rxctrlout       : out    vl_logic_vector(3 downto 0);
        rxdataout       : out    vl_logic_vector(31 downto 0);
        rxdigitalresetout: out    vl_logic_vector(3 downto 0);
        rxibpowerdown   : out    vl_logic_vector(3 downto 0);
        rxphfifox4byteselout: out    vl_logic;
        rxphfifox4rdenableout: out    vl_logic;
        rxphfifox4wrclkout: out    vl_logic;
        rxphfifox4wrenableout: out    vl_logic;
        testout         : out    vl_logic_vector(2399 downto 0);
        txanalogresetout: out    vl_logic_vector(3 downto 0);
        txctrlout       : out    vl_logic_vector(3 downto 0);
        txdataout       : out    vl_logic_vector(31 downto 0);
        txdetectrxpowerdown: out    vl_logic_vector(3 downto 0);
        txdigitalresetout: out    vl_logic_vector(3 downto 0);
        txdividerpowerdown: out    vl_logic_vector(3 downto 0);
        txobpowerdown   : out    vl_logic_vector(3 downto 0);
        txphfifox4byteselout: out    vl_logic;
        txphfifox4rdclkout: out    vl_logic;
        txphfifox4rdenableout: out    vl_logic;
        txphfifox4wrenableout: out    vl_logic;
        rxpmadprioout   : out    vl_logic_vector(1199 downto 0);
        rxpcsdprioout   : out    vl_logic_vector(1599 downto 0);
        txpmadprioout   : out    vl_logic_vector(1199 downto 0);
        txpcsdprioout   : out    vl_logic_vector(599 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of auto_spd_deassert_ph_fifo_rst_count : constant is 1;
    attribute mti_svvh_generic_type of auto_spd_phystatus_notify_count : constant is 1;
    attribute mti_svvh_generic_type of coreclk_out_gated_by_quad_reset : constant is 1;
    attribute mti_svvh_generic_type of in_xaui_mode : constant is 1;
    attribute mti_svvh_generic_type of pipe_auto_speed_nego_enable : constant is 1;
    attribute mti_svvh_generic_type of rx_xaui_sm_backward_compatible_enable : constant is 1;
    attribute mti_svvh_generic_type of rx0_channel_bonding : constant is 1;
    attribute mti_svvh_generic_type of rx0_clk1_mux_select : constant is 1;
    attribute mti_svvh_generic_type of rx0_clk2_mux_select : constant is 1;
    attribute mti_svvh_generic_type of rx0_clk_pd_enable : constant is 1;
    attribute mti_svvh_generic_type of rx0_ph_fifo_reg_mode : constant is 1;
    attribute mti_svvh_generic_type of rx0_ph_fifo_reset_enable : constant is 1;
    attribute mti_svvh_generic_type of rx0_ph_fifo_user_ctrl_enable : constant is 1;
    attribute mti_svvh_generic_type of rx0_rd_clk_mux_select : constant is 1;
    attribute mti_svvh_generic_type of rx0_recovered_clk_mux_select : constant is 1;
    attribute mti_svvh_generic_type of rx0_reset_clock_output_during_digital_reset : constant is 1;
    attribute mti_svvh_generic_type of rx0_use_double_data_mode : constant is 1;
    attribute mti_svvh_generic_type of select_refclk_dig : constant is 1;
    attribute mti_svvh_generic_type of tx_xaui_sm_backward_compatible_enable : constant is 1;
    attribute mti_svvh_generic_type of tx0_channel_bonding : constant is 1;
    attribute mti_svvh_generic_type of tx0_clk_pd_enable : constant is 1;
    attribute mti_svvh_generic_type of tx0_ph_fifo_reset_enable : constant is 1;
    attribute mti_svvh_generic_type of tx0_ph_fifo_user_ctrl_enable : constant is 1;
    attribute mti_svvh_generic_type of tx0_rd_clk_mux_select : constant is 1;
    attribute mti_svvh_generic_type of tx0_reset_clock_output_during_digital_reset : constant is 1;
    attribute mti_svvh_generic_type of tx0_use_double_data_mode : constant is 1;
    attribute mti_svvh_generic_type of tx0_wr_clk_mux_select : constant is 1;
    attribute mti_svvh_generic_type of use_coreclk_out_post_divider : constant is 1;
    attribute mti_svvh_generic_type of use_deskew_fifo : constant is 1;
    attribute mti_svvh_generic_type of dprio_config_mode : constant is 1;
    attribute mti_svvh_generic_type of rx_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of tx_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of pll_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of portaddr : constant is 1;
    attribute mti_svvh_generic_type of devaddr : constant is 1;
    attribute mti_svvh_generic_type of rx0_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of rx1_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of rx2_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of rx3_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of tx0_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of tx1_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of tx2_logical_to_physical_mapping : constant is 1;
    attribute mti_svvh_generic_type of tx3_logical_to_physical_mapping : constant is 1;
end cycloneiv_hssi_cmu;
