library verilog;
use verilog.vl_types.all;
entity cycloneiv_hssi_cmu_dprio_centrl_bus_out_mux is
    port(
        centrl_ctrl_in1 : in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in2 : in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in3 : in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in4 : in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in5 : in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in6 : in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in7 : in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in8 : in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in9 : in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in10: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in11: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in12: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in13: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in14: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in15: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in16: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in17: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in18: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in19: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in20: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in21: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in22: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in23: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in24: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in25: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in26: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in27: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in28: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in29: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in30: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in31: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in32: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in33: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in34: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in35: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in36: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in37: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in38: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in39: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in40: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in41: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in42: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in43: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in44: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in45: in     vl_logic_vector(15 downto 0);
        centrl_ctrl_in46: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in1: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in2: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in3: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in4: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in5: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in6: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in7: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in8: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in9: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in10: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in11: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in12: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in13: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in14: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in15: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in16: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in17: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in18: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in19: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in20: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in21: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in22: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in23: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in24: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in25: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in26: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in27: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in28: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in29: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in30: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in31: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in32: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in33: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in34: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in35: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in36: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in37: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in38: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in39: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in40: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in41: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in42: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in43: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in44: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in45: in     vl_logic_vector(15 downto 0);
        hw_address_ctrl_in46: in     vl_logic_vector(15 downto 0);
        reg_addr        : in     vl_logic_vector(15 downto 0);
        centrl_ctrl_out : out    vl_logic_vector(15 downto 0)
    );
end cycloneiv_hssi_cmu_dprio_centrl_bus_out_mux;
