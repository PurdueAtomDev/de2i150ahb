library verilog;
use verilog.vl_types.all;
entity test_program is
end test_program;
