library verilog;
use verilog.vl_types.all;
entity cycloneiv_hssi_rx_pma is
    generic(
        lpm_type        : string  := "cycloneiv_hssi_rx_pma";
        allow_serial_loopback: string  := "false";
        channel_number  : integer := 0;
        common_mode     : string  := "0.82V";
        deserialization_factor: integer := 8;
        dprio_config_mode: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        enable_local_divider: string  := "false";
        enable_dpa_shift: string  := "false";
        enable_initial_phase_selection: string  := "false";
        enable_pd_counter_accumulate_mode: string  := "false";
        enable_ltd      : string  := "false";
        enable_ltr      : string  := "false";
        eq_dc_gain      : integer := 0;
        eq_setting      : integer := 1;
        force_signal_detect: string  := "true";
        initial_phase_value: integer := 0;
        logical_channel_address: integer := 0;
        offset_cancellation: integer := 0;
        pd1_counter_setting: integer := 5;
        pd2_counter_setting: integer := 5;
        pd_rising_edge_only: string  := "false";
        phase_step_add_setting: integer := 2;
        phase_step_sub_setting: integer := 1;
        pi_frequency_selector: integer := 0;
        ppm_gen1_2_xcnt_en: integer := 1;
        ppm_post_eidle  : integer := 0;
        ppmselect       : integer := 0;
        protocol_hint   : string  := "basic";
        effective_data_rate: string  := "unused";
        send_reverse_serial_loopback_data: string  := "false";
        send_reverse_serial_loopback_recovered_clk: string  := "false";
        signal_detect_hysteresis: integer := 4;
        signal_detect_hysteresis_valid_threshold: integer := 1;
        signal_detect_loss_threshold: integer := 1;
        termination     : string  := "OCT 100 Ohms";
        use_external_termination: string  := "false";
        loop_1_digital_filter: integer := 8;
        enable_second_order_loop: string  := "false"
    );
    port(
        crupowerdn      : in     vl_logic;
        datain          : in     vl_logic;
        deserclock      : in     vl_logic;
        dpashift        : in     vl_logic;
        dpriodisable    : in     vl_logic;
        dprioin         : in     vl_logic_vector(299 downto 0);
        locktodata      : in     vl_logic;
        locktoref       : in     vl_logic;
        powerdn         : in     vl_logic;
        ppmdetectrefclk : in     vl_logic;
        rxpmareset      : in     vl_logic;
        seriallpbkin    : in     vl_logic;
        testbussel      : in     vl_logic_vector(3 downto 0);
        analogtestbus   : out    vl_logic_vector(7 downto 0);
        clockout        : out    vl_logic;
        datastrobeout   : out    vl_logic;
        dprioout        : out    vl_logic_vector(299 downto 0);
        diagnosticlpbkout: out    vl_logic;
        freqlocked      : out    vl_logic;
        locktorefout    : out    vl_logic;
        recoverdataout  : out    vl_logic_vector(9 downto 0);
        reverselpbkout  : out    vl_logic;
        signaldetect    : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of allow_serial_loopback : constant is 1;
    attribute mti_svvh_generic_type of channel_number : constant is 1;
    attribute mti_svvh_generic_type of common_mode : constant is 1;
    attribute mti_svvh_generic_type of deserialization_factor : constant is 1;
    attribute mti_svvh_generic_type of dprio_config_mode : constant is 1;
    attribute mti_svvh_generic_type of enable_local_divider : constant is 1;
    attribute mti_svvh_generic_type of enable_dpa_shift : constant is 1;
    attribute mti_svvh_generic_type of enable_initial_phase_selection : constant is 1;
    attribute mti_svvh_generic_type of enable_pd_counter_accumulate_mode : constant is 1;
    attribute mti_svvh_generic_type of enable_ltd : constant is 1;
    attribute mti_svvh_generic_type of enable_ltr : constant is 1;
    attribute mti_svvh_generic_type of eq_dc_gain : constant is 1;
    attribute mti_svvh_generic_type of eq_setting : constant is 1;
    attribute mti_svvh_generic_type of force_signal_detect : constant is 1;
    attribute mti_svvh_generic_type of initial_phase_value : constant is 1;
    attribute mti_svvh_generic_type of logical_channel_address : constant is 1;
    attribute mti_svvh_generic_type of offset_cancellation : constant is 1;
    attribute mti_svvh_generic_type of pd1_counter_setting : constant is 1;
    attribute mti_svvh_generic_type of pd2_counter_setting : constant is 1;
    attribute mti_svvh_generic_type of pd_rising_edge_only : constant is 1;
    attribute mti_svvh_generic_type of phase_step_add_setting : constant is 1;
    attribute mti_svvh_generic_type of phase_step_sub_setting : constant is 1;
    attribute mti_svvh_generic_type of pi_frequency_selector : constant is 1;
    attribute mti_svvh_generic_type of ppm_gen1_2_xcnt_en : constant is 1;
    attribute mti_svvh_generic_type of ppm_post_eidle : constant is 1;
    attribute mti_svvh_generic_type of ppmselect : constant is 1;
    attribute mti_svvh_generic_type of protocol_hint : constant is 1;
    attribute mti_svvh_generic_type of effective_data_rate : constant is 1;
    attribute mti_svvh_generic_type of send_reverse_serial_loopback_data : constant is 1;
    attribute mti_svvh_generic_type of send_reverse_serial_loopback_recovered_clk : constant is 1;
    attribute mti_svvh_generic_type of signal_detect_hysteresis : constant is 1;
    attribute mti_svvh_generic_type of signal_detect_hysteresis_valid_threshold : constant is 1;
    attribute mti_svvh_generic_type of signal_detect_loss_threshold : constant is 1;
    attribute mti_svvh_generic_type of termination : constant is 1;
    attribute mti_svvh_generic_type of use_external_termination : constant is 1;
    attribute mti_svvh_generic_type of loop_1_digital_filter : constant is 1;
    attribute mti_svvh_generic_type of enable_second_order_loop : constant is 1;
end cycloneiv_hssi_rx_pma;
