library verilog;
use verilog.vl_types.all;
entity cycloneiv_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end cycloneiv_routing_wire;
