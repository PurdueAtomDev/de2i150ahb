library verilog;
use verilog.vl_types.all;
entity avalon_utilities_pkg is
end avalon_utilities_pkg;
