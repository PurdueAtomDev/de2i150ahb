// ahb_master_slave_with_pcie.v

// Generated using ACDS version 14.0 200 at 2015.08.10.15:09:47

`timescale 1 ps / 1 ps
module ahb_master_slave_with_pcie (
		input  wire        clk_clk,                                       //                              clk.clk
		input  wire        reset_reset_n,                                 //                            reset.reset_n
		input  wire [3:0]  pcie_ip_reconfig_togxb_data,                   //           pcie_ip_reconfig_togxb.data
		input  wire        pcie_ip_refclk_export,                         //                   pcie_ip_refclk.export
		input  wire [39:0] pcie_ip_test_in_test_in,                       //                  pcie_ip_test_in.test_in
		input  wire        pcie_ip_pcie_rstn_export,                      //                pcie_ip_pcie_rstn.export
		output wire        pcie_ip_clocks_sim_clk250_export,              //               pcie_ip_clocks_sim.clk250_export
		output wire        pcie_ip_clocks_sim_clk500_export,              //                                 .clk500_export
		output wire        pcie_ip_clocks_sim_clk125_export,              //                                 .clk125_export
		input  wire        pcie_ip_reconfig_busy_busy_altgxb_reconfig,    //            pcie_ip_reconfig_busy.busy_altgxb_reconfig
		input  wire        pcie_ip_pipe_ext_pipe_mode,                    //                 pcie_ip_pipe_ext.pipe_mode
		input  wire        pcie_ip_pipe_ext_phystatus_ext,                //                                 .phystatus_ext
		output wire        pcie_ip_pipe_ext_rate_ext,                     //                                 .rate_ext
		output wire [1:0]  pcie_ip_pipe_ext_powerdown_ext,                //                                 .powerdown_ext
		output wire        pcie_ip_pipe_ext_txdetectrx_ext,               //                                 .txdetectrx_ext
		input  wire        pcie_ip_pipe_ext_rxelecidle0_ext,              //                                 .rxelecidle0_ext
		input  wire [7:0]  pcie_ip_pipe_ext_rxdata0_ext,                  //                                 .rxdata0_ext
		input  wire [2:0]  pcie_ip_pipe_ext_rxstatus0_ext,                //                                 .rxstatus0_ext
		input  wire        pcie_ip_pipe_ext_rxvalid0_ext,                 //                                 .rxvalid0_ext
		input  wire        pcie_ip_pipe_ext_rxdatak0_ext,                 //                                 .rxdatak0_ext
		output wire [7:0]  pcie_ip_pipe_ext_txdata0_ext,                  //                                 .txdata0_ext
		output wire        pcie_ip_pipe_ext_txdatak0_ext,                 //                                 .txdatak0_ext
		output wire        pcie_ip_pipe_ext_rxpolarity0_ext,              //                                 .rxpolarity0_ext
		output wire        pcie_ip_pipe_ext_txcompl0_ext,                 //                                 .txcompl0_ext
		output wire        pcie_ip_pipe_ext_txelecidle0_ext,              //                                 .txelecidle0_ext
		input  wire        pcie_ip_rx_in_rx_datain_0,                     //                    pcie_ip_rx_in.rx_datain_0
		output wire        pcie_ip_tx_out_tx_dataout_0,                   //                   pcie_ip_tx_out.tx_dataout_0
		output wire [4:0]  pcie_ip_reconfig_fromgxb_0_data,               //       pcie_ip_reconfig_fromgxb_0.data
		output wire [11:0] sdram_addr,                                    //                            sdram.addr
		output wire [1:0]  sdram_ba,                                      //                                 .ba
		output wire        sdram_cas_n,                                   //                                 .cas_n
		output wire        sdram_cke,                                     //                                 .cke
		output wire        sdram_cs_n,                                    //                                 .cs_n
		inout  wire [31:0] sdram_dq,                                      //                                 .dq
		output wire [3:0]  sdram_dqm,                                     //                                 .dqm
		output wire        sdram_ras_n,                                   //                                 .ras_n
		output wire        sdram_we_n,                                    //                                 .we_n
		output wire        altpll_sdram_clk,                              //                     altpll_sdram.clk
		input  wire        pcie_ip_powerdown_pll_powerdown,               //                pcie_ip_powerdown.pll_powerdown
		input  wire        pcie_ip_powerdown_gxb_powerdown,               //                                 .gxb_powerdown
		input  wire        ahb_master_slave_2_0_conduit_end_add_data_sel, // ahb_master_slave_2_0_conduit_end.add_data_sel
		input  wire [15:0] ahb_master_slave_2_0_conduit_end_rdwr_address, //                                 .rdwr_address
		output wire [31:0] ahb_master_slave_2_0_conduit_end_display_data  //                                 .display_data
	);

	wire         pcie_ip_pcie_core_clk_clk;                                        // pcie_ip:pcie_core_clk_clk -> [irq_mapper:clk, mm_interconnect_0:pcie_ip_pcie_core_clk_clk, mm_interconnect_1:pcie_ip_pcie_core_clk_clk, mm_interconnect_2:pcie_ip_pcie_core_clk_clk, pcie_ip:fixedclk_clk, rst_controller:clk, rst_controller_003:clk, sgdma:clk]
	wire         altpll_qsys_c3_clk;                                               // altpll_qsys:c3 -> [pcie_ip:cal_blk_clk_clk, pcie_ip:reconfig_gxbclk_clk]
	wire         avalon2ahb_bridge_0_ahb_master_hwrite;                            // avalon2ahb_bridge_0:HWRITE -> ahb_master_slave_2_0:slave_HWRITE
	wire  [31:0] avalon2ahb_bridge_0_ahb_master_hwdata;                            // avalon2ahb_bridge_0:HWDATA -> ahb_master_slave_2_0:slave_HWDATA
	wire   [3:0] avalon2ahb_bridge_0_ahb_master_hprot;                             // avalon2ahb_bridge_0:HPROT -> ahb_master_slave_2_0:slave_HPROT
	wire         avalon2ahb_bridge_0_ahb_master_hreadyin;                          // avalon2ahb_bridge_0:HREADYIN -> ahb_master_slave_2_0:slave_HREADY
	wire   [2:0] avalon2ahb_bridge_0_ahb_master_hsize;                             // avalon2ahb_bridge_0:HSIZE -> ahb_master_slave_2_0:slave_HSIZE
	wire  [31:0] avalon2ahb_bridge_0_ahb_master_hrdata;                            // ahb_master_slave_2_0:slave_HRDATA -> avalon2ahb_bridge_0:HRDATA
	wire         avalon2ahb_bridge_0_ahb_master_hsel;                              // avalon2ahb_bridge_0:HSEL -> ahb_master_slave_2_0:slave_HSEL
	wire   [1:0] avalon2ahb_bridge_0_ahb_master_htrans;                            // avalon2ahb_bridge_0:HTRANS -> ahb_master_slave_2_0:slave_HTRANS
	wire   [1:0] avalon2ahb_bridge_0_ahb_master_hresp;                             // ahb_master_slave_2_0:slave_HRESP -> avalon2ahb_bridge_0:HRESP
	wire  [31:0] avalon2ahb_bridge_0_ahb_master_haddr;                             // avalon2ahb_bridge_0:HADDR -> ahb_master_slave_2_0:slave_HADDR
	wire         avalon2ahb_bridge_0_ahb_master_hready;                            // ahb_master_slave_2_0:slave_HREADYOUT -> avalon2ahb_bridge_0:HREADY
	wire   [2:0] avalon2ahb_bridge_0_ahb_master_hburst;                            // avalon2ahb_bridge_0:HBURST -> ahb_master_slave_2_0:slave_HBURST
	wire         ahb_master_slave_2_0_ahb_master_hwrite;                           // ahb_master_slave_2_0:master_HWRITE -> ahb2avalon_burst_bridge_0:HWRITE
	wire  [31:0] ahb_master_slave_2_0_ahb_master_hwdata;                           // ahb_master_slave_2_0:master_HWDATA -> ahb2avalon_burst_bridge_0:HWDATA
	wire   [3:0] ahb_master_slave_2_0_ahb_master_hprot;                            // ahb_master_slave_2_0:master_HPROT -> ahb2avalon_burst_bridge_0:HPROT
	wire         ahb_master_slave_2_0_ahb_master_hreadyin;                         // ahb_master_slave_2_0:master_HREADYIN -> ahb2avalon_burst_bridge_0:HREADY
	wire   [2:0] ahb_master_slave_2_0_ahb_master_hsize;                            // ahb_master_slave_2_0:master_HSIZE -> ahb2avalon_burst_bridge_0:HSIZE
	wire  [31:0] ahb_master_slave_2_0_ahb_master_hrdata;                           // ahb2avalon_burst_bridge_0:HRDATA -> ahb_master_slave_2_0:master_HRDATA
	wire         ahb_master_slave_2_0_ahb_master_hsel;                             // ahb_master_slave_2_0:master_HSEL -> ahb2avalon_burst_bridge_0:HSEL
	wire   [1:0] ahb_master_slave_2_0_ahb_master_htrans;                           // ahb_master_slave_2_0:master_HTRANS -> ahb2avalon_burst_bridge_0:HTRANS
	wire   [1:0] ahb_master_slave_2_0_ahb_master_hresp;                            // ahb2avalon_burst_bridge_0:HRESP -> ahb_master_slave_2_0:master_HRESP
	wire         ahb_master_slave_2_0_ahb_master_hready;                           // ahb2avalon_burst_bridge_0:HREADYOUT -> ahb_master_slave_2_0:master_HREADY
	wire  [31:0] ahb_master_slave_2_0_ahb_master_haddr;                            // ahb_master_slave_2_0:master_HADDR -> ahb2avalon_burst_bridge_0:HADDR
	wire   [2:0] ahb_master_slave_2_0_ahb_master_hburst;                           // ahb_master_slave_2_0:master_HBURST -> ahb2avalon_burst_bridge_0:HBURST
	wire   [6:0] pcie_ip_bar2_burstcount;                                          // pcie_ip:bar2_burstcount -> mm_interconnect_0:pcie_ip_bar2_burstcount
	wire         pcie_ip_bar2_waitrequest;                                         // mm_interconnect_0:pcie_ip_bar2_waitrequest -> pcie_ip:bar2_waitrequest
	wire  [63:0] pcie_ip_bar2_writedata;                                           // pcie_ip:bar2_writedata -> mm_interconnect_0:pcie_ip_bar2_writedata
	wire  [31:0] pcie_ip_bar2_address;                                             // pcie_ip:bar2_address -> mm_interconnect_0:pcie_ip_bar2_address
	wire         pcie_ip_bar2_write;                                               // pcie_ip:bar2_write -> mm_interconnect_0:pcie_ip_bar2_write
	wire         pcie_ip_bar2_read;                                                // pcie_ip:bar2_read -> mm_interconnect_0:pcie_ip_bar2_read
	wire  [63:0] pcie_ip_bar2_readdata;                                            // mm_interconnect_0:pcie_ip_bar2_readdata -> pcie_ip:bar2_readdata
	wire   [7:0] pcie_ip_bar2_byteenable;                                          // pcie_ip:bar2_byteenable -> mm_interconnect_0:pcie_ip_bar2_byteenable
	wire         pcie_ip_bar2_readdatavalid;                                       // mm_interconnect_0:pcie_ip_bar2_readdatavalid -> pcie_ip:bar2_readdatavalid
	wire  [31:0] mm_interconnect_0_sgdma_csr_writedata;                            // mm_interconnect_0:sgdma_csr_writedata -> sgdma:csr_writedata
	wire   [3:0] mm_interconnect_0_sgdma_csr_address;                              // mm_interconnect_0:sgdma_csr_address -> sgdma:csr_address
	wire         mm_interconnect_0_sgdma_csr_chipselect;                           // mm_interconnect_0:sgdma_csr_chipselect -> sgdma:csr_chipselect
	wire         mm_interconnect_0_sgdma_csr_write;                                // mm_interconnect_0:sgdma_csr_write -> sgdma:csr_write
	wire         mm_interconnect_0_sgdma_csr_read;                                 // mm_interconnect_0:sgdma_csr_read -> sgdma:csr_read
	wire  [31:0] mm_interconnect_0_sgdma_csr_readdata;                             // sgdma:csr_readdata -> mm_interconnect_0:sgdma_csr_readdata
	wire         mm_interconnect_0_pcie_ip_cra_waitrequest;                        // pcie_ip:cra_waitrequest -> mm_interconnect_0:pcie_ip_cra_waitrequest
	wire  [31:0] mm_interconnect_0_pcie_ip_cra_writedata;                          // mm_interconnect_0:pcie_ip_cra_writedata -> pcie_ip:cra_writedata
	wire  [11:0] mm_interconnect_0_pcie_ip_cra_address;                            // mm_interconnect_0:pcie_ip_cra_address -> pcie_ip:cra_address
	wire         mm_interconnect_0_pcie_ip_cra_chipselect;                         // mm_interconnect_0:pcie_ip_cra_chipselect -> pcie_ip:cra_chipselect
	wire         mm_interconnect_0_pcie_ip_cra_write;                              // mm_interconnect_0:pcie_ip_cra_write -> pcie_ip:cra_write
	wire         mm_interconnect_0_pcie_ip_cra_read;                               // mm_interconnect_0:pcie_ip_cra_read -> pcie_ip:cra_read
	wire  [31:0] mm_interconnect_0_pcie_ip_cra_readdata;                           // pcie_ip:cra_readdata -> mm_interconnect_0:pcie_ip_cra_readdata
	wire   [3:0] mm_interconnect_0_pcie_ip_cra_byteenable;                         // mm_interconnect_0:pcie_ip_cra_byteenable -> pcie_ip:cra_byteenable
	wire         sgdma_descriptor_read_waitrequest;                                // mm_interconnect_1:sgdma_descriptor_read_waitrequest -> sgdma:descriptor_read_waitrequest
	wire  [31:0] sgdma_descriptor_read_address;                                    // sgdma:descriptor_read_address -> mm_interconnect_1:sgdma_descriptor_read_address
	wire         sgdma_descriptor_read_read;                                       // sgdma:descriptor_read_read -> mm_interconnect_1:sgdma_descriptor_read_read
	wire  [31:0] sgdma_descriptor_read_readdata;                                   // mm_interconnect_1:sgdma_descriptor_read_readdata -> sgdma:descriptor_read_readdata
	wire         sgdma_descriptor_read_readdatavalid;                              // mm_interconnect_1:sgdma_descriptor_read_readdatavalid -> sgdma:descriptor_read_readdatavalid
	wire         sgdma_descriptor_write_waitrequest;                               // mm_interconnect_1:sgdma_descriptor_write_waitrequest -> sgdma:descriptor_write_waitrequest
	wire  [31:0] sgdma_descriptor_write_writedata;                                 // sgdma:descriptor_write_writedata -> mm_interconnect_1:sgdma_descriptor_write_writedata
	wire  [31:0] sgdma_descriptor_write_address;                                   // sgdma:descriptor_write_address -> mm_interconnect_1:sgdma_descriptor_write_address
	wire         sgdma_descriptor_write_write;                                     // sgdma:descriptor_write_write -> mm_interconnect_1:sgdma_descriptor_write_write
	wire   [3:0] sgdma_m_read_burstcount;                                          // sgdma:m_read_burstcount -> mm_interconnect_1:sgdma_m_read_burstcount
	wire         sgdma_m_read_waitrequest;                                         // mm_interconnect_1:sgdma_m_read_waitrequest -> sgdma:m_read_waitrequest
	wire  [31:0] sgdma_m_read_address;                                             // sgdma:m_read_address -> mm_interconnect_1:sgdma_m_read_address
	wire         sgdma_m_read_read;                                                // sgdma:m_read_read -> mm_interconnect_1:sgdma_m_read_read
	wire  [31:0] sgdma_m_read_readdata;                                            // mm_interconnect_1:sgdma_m_read_readdata -> sgdma:m_read_readdata
	wire         sgdma_m_read_readdatavalid;                                       // mm_interconnect_1:sgdma_m_read_readdatavalid -> sgdma:m_read_readdatavalid
	wire   [7:0] sgdma_m_write_burstcount;                                         // sgdma:m_write_burstcount -> mm_interconnect_1:sgdma_m_write_burstcount
	wire         sgdma_m_write_waitrequest;                                        // mm_interconnect_1:sgdma_m_write_waitrequest -> sgdma:m_write_waitrequest
	wire  [31:0] sgdma_m_write_writedata;                                          // sgdma:m_write_writedata -> mm_interconnect_1:sgdma_m_write_writedata
	wire  [31:0] sgdma_m_write_address;                                            // sgdma:m_write_address -> mm_interconnect_1:sgdma_m_write_address
	wire         sgdma_m_write_write;                                              // sgdma:m_write_write -> mm_interconnect_1:sgdma_m_write_write
	wire   [3:0] sgdma_m_write_byteenable;                                         // sgdma:m_write_byteenable -> mm_interconnect_1:sgdma_m_write_byteenable
	wire   [3:0] ahb2avalon_burst_bridge_0_avalon_master_burstcount;               // ahb2avalon_burst_bridge_0:burstcount -> mm_interconnect_1:ahb2avalon_burst_bridge_0_avalon_master_burstcount
	wire         ahb2avalon_burst_bridge_0_avalon_master_waitrequest;              // mm_interconnect_1:ahb2avalon_burst_bridge_0_avalon_master_waitrequest -> ahb2avalon_burst_bridge_0:waitrequest
	wire  [31:0] ahb2avalon_burst_bridge_0_avalon_master_writedata;                // ahb2avalon_burst_bridge_0:writedata -> mm_interconnect_1:ahb2avalon_burst_bridge_0_avalon_master_writedata
	wire  [31:0] ahb2avalon_burst_bridge_0_avalon_master_address;                  // ahb2avalon_burst_bridge_0:address -> mm_interconnect_1:ahb2avalon_burst_bridge_0_avalon_master_address
	wire         ahb2avalon_burst_bridge_0_avalon_master_write;                    // ahb2avalon_burst_bridge_0:write -> mm_interconnect_1:ahb2avalon_burst_bridge_0_avalon_master_write
	wire         ahb2avalon_burst_bridge_0_avalon_master_read;                     // ahb2avalon_burst_bridge_0:read -> mm_interconnect_1:ahb2avalon_burst_bridge_0_avalon_master_read
	wire  [31:0] ahb2avalon_burst_bridge_0_avalon_master_readdata;                 // mm_interconnect_1:ahb2avalon_burst_bridge_0_avalon_master_readdata -> ahb2avalon_burst_bridge_0:readdata
	wire         ahb2avalon_burst_bridge_0_avalon_master_readdatavalid;            // mm_interconnect_1:ahb2avalon_burst_bridge_0_avalon_master_readdatavalid -> ahb2avalon_burst_bridge_0:readdatavalid
	wire   [3:0] ahb2avalon_burst_bridge_0_avalon_master_byteenable;               // ahb2avalon_burst_bridge_0:byteenable -> mm_interconnect_1:ahb2avalon_burst_bridge_0_avalon_master_byteenable
	wire         mm_interconnect_1_pcie_ip_txs_waitrequest;                        // pcie_ip:txs_waitrequest -> mm_interconnect_1:pcie_ip_txs_waitrequest
	wire   [6:0] mm_interconnect_1_pcie_ip_txs_burstcount;                         // mm_interconnect_1:pcie_ip_txs_burstcount -> pcie_ip:txs_burstcount
	wire  [63:0] mm_interconnect_1_pcie_ip_txs_writedata;                          // mm_interconnect_1:pcie_ip_txs_writedata -> pcie_ip:txs_writedata
	wire  [30:0] mm_interconnect_1_pcie_ip_txs_address;                            // mm_interconnect_1:pcie_ip_txs_address -> pcie_ip:txs_address
	wire         mm_interconnect_1_pcie_ip_txs_chipselect;                         // mm_interconnect_1:pcie_ip_txs_chipselect -> pcie_ip:txs_chipselect
	wire         mm_interconnect_1_pcie_ip_txs_write;                              // mm_interconnect_1:pcie_ip_txs_write -> pcie_ip:txs_write
	wire         mm_interconnect_1_pcie_ip_txs_read;                               // mm_interconnect_1:pcie_ip_txs_read -> pcie_ip:txs_read
	wire  [63:0] mm_interconnect_1_pcie_ip_txs_readdata;                           // pcie_ip:txs_readdata -> mm_interconnect_1:pcie_ip_txs_readdata
	wire         mm_interconnect_1_pcie_ip_txs_readdatavalid;                      // pcie_ip:txs_readdatavalid -> mm_interconnect_1:pcie_ip_txs_readdatavalid
	wire   [7:0] mm_interconnect_1_pcie_ip_txs_byteenable;                         // mm_interconnect_1:pcie_ip_txs_byteenable -> pcie_ip:txs_byteenable
	wire         mm_interconnect_1_sdram_s1_waitrequest;                           // sdram:za_waitrequest -> mm_interconnect_1:sdram_s1_waitrequest
	wire  [31:0] mm_interconnect_1_sdram_s1_writedata;                             // mm_interconnect_1:sdram_s1_writedata -> sdram:az_data
	wire  [23:0] mm_interconnect_1_sdram_s1_address;                               // mm_interconnect_1:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_1_sdram_s1_chipselect;                            // mm_interconnect_1:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_1_sdram_s1_write;                                 // mm_interconnect_1:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_1_sdram_s1_read;                                  // mm_interconnect_1:sdram_s1_read -> sdram:az_rd_n
	wire  [31:0] mm_interconnect_1_sdram_s1_readdata;                              // sdram:za_data -> mm_interconnect_1:sdram_s1_readdata
	wire         mm_interconnect_1_sdram_s1_readdatavalid;                         // sdram:za_valid -> mm_interconnect_1:sdram_s1_readdatavalid
	wire   [3:0] mm_interconnect_1_sdram_s1_byteenable;                            // mm_interconnect_1:sdram_s1_byteenable -> sdram:az_be_n
	wire   [6:0] pcie_ip_bar1_0_burstcount;                                        // pcie_ip:bar1_0_burstcount -> mm_interconnect_2:pcie_ip_bar1_0_burstcount
	wire         pcie_ip_bar1_0_waitrequest;                                       // mm_interconnect_2:pcie_ip_bar1_0_waitrequest -> pcie_ip:bar1_0_waitrequest
	wire  [63:0] pcie_ip_bar1_0_writedata;                                         // pcie_ip:bar1_0_writedata -> mm_interconnect_2:pcie_ip_bar1_0_writedata
	wire  [31:0] pcie_ip_bar1_0_address;                                           // pcie_ip:bar1_0_address -> mm_interconnect_2:pcie_ip_bar1_0_address
	wire         pcie_ip_bar1_0_write;                                             // pcie_ip:bar1_0_write -> mm_interconnect_2:pcie_ip_bar1_0_write
	wire         pcie_ip_bar1_0_read;                                              // pcie_ip:bar1_0_read -> mm_interconnect_2:pcie_ip_bar1_0_read
	wire  [63:0] pcie_ip_bar1_0_readdata;                                          // mm_interconnect_2:pcie_ip_bar1_0_readdata -> pcie_ip:bar1_0_readdata
	wire   [7:0] pcie_ip_bar1_0_byteenable;                                        // pcie_ip:bar1_0_byteenable -> mm_interconnect_2:pcie_ip_bar1_0_byteenable
	wire         pcie_ip_bar1_0_readdatavalid;                                     // mm_interconnect_2:pcie_ip_bar1_0_readdatavalid -> pcie_ip:bar1_0_readdatavalid
	wire         mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_waitrequest;   // avalon2ahb_bridge_0:waitrequest -> mm_interconnect_2:avalon2ahb_bridge_0_avalon_slave_waitrequest
	wire  [31:0] mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_writedata;     // mm_interconnect_2:avalon2ahb_bridge_0_avalon_slave_writedata -> avalon2ahb_bridge_0:writedata
	wire   [4:0] mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_address;       // mm_interconnect_2:avalon2ahb_bridge_0_avalon_slave_address -> avalon2ahb_bridge_0:address
	wire         mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_write;         // mm_interconnect_2:avalon2ahb_bridge_0_avalon_slave_write -> avalon2ahb_bridge_0:write
	wire         mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_read;          // mm_interconnect_2:avalon2ahb_bridge_0_avalon_slave_read -> avalon2ahb_bridge_0:read
	wire  [31:0] mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_readdata;      // avalon2ahb_bridge_0:readdata -> mm_interconnect_2:avalon2ahb_bridge_0_avalon_slave_readdata
	wire         mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_readdatavalid; // avalon2ahb_bridge_0:readdatavalid -> mm_interconnect_2:avalon2ahb_bridge_0_avalon_slave_readdatavalid
	wire         irq_mapper_receiver0_irq;                                         // sgdma:csr_irq -> irq_mapper:receiver0_irq
	wire  [15:0] pcie_ip_rxm_irq_irq;                                              // irq_mapper:sender_irq -> pcie_ip:rxm_irq_irq
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [mm_interconnect_0:sgdma_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sgdma_reset_reset_bridge_in_reset_reset, sgdma:system_reset_n]
	wire         pcie_ip_pcie_core_reset_reset;                                    // pcie_ip:pcie_core_reset_reset_n -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_003:reset_in0]
	wire         rst_controller_001_reset_out_reset;                               // rst_controller_001:reset_out -> [altpll_qsys:reset, mm_interconnect_1:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]
	wire         rst_controller_002_reset_out_reset;                               // rst_controller_002:reset_out -> [ahb2avalon_burst_bridge_0:reset_n, ahb_master_slave_2_0:HRESETn, avalon2ahb_bridge_0:reset_n, mm_interconnect_1:ahb2avalon_burst_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:avalon2ahb_bridge_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_003_reset_out_reset;                               // rst_controller_003:reset_out -> [irq_mapper:reset, mm_interconnect_0:pcie_ip_bar2_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pcie_ip_txs_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset_reset]

	ahb_master_slave_with_pcie_pcie_ip #(
		.p_pcie_hip_type                     ("2"),
		.lane_mask                           (8'b11111110),
		.max_link_width                      (1),
		.millisecond_cycle_count             ("125000"),
		.enable_gen2_core                    ("false"),
		.gen2_lane_rate_mode                 ("false"),
		.no_soft_reset                       ("false"),
		.core_clk_divider                    (2),
		.enable_ch0_pclk_out                 ("true"),
		.core_clk_source                     ("pclk"),
		.CB_P2A_AVALON_ADDR_B0               (0),
		.bar0_size_mask                      (7),
		.bar0_io_space                       ("false"),
		.bar0_64bit_mem_space                ("true"),
		.bar0_prefetchable                   ("true"),
		.CB_P2A_AVALON_ADDR_B1               (0),
		.bar1_size_mask                      (0),
		.bar1_io_space                       ("false"),
		.bar1_64bit_mem_space                ("true"),
		.bar1_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B2               (0),
		.bar2_size_mask                      (15),
		.bar2_io_space                       ("false"),
		.bar2_64bit_mem_space                ("false"),
		.bar2_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B3               (0),
		.bar3_size_mask                      (0),
		.bar3_io_space                       ("false"),
		.bar3_64bit_mem_space                ("false"),
		.bar3_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B4               (0),
		.bar4_size_mask                      (0),
		.bar4_io_space                       ("false"),
		.bar4_64bit_mem_space                ("false"),
		.bar4_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B5               (0),
		.bar5_size_mask                      (0),
		.bar5_io_space                       ("false"),
		.bar5_64bit_mem_space                ("false"),
		.bar5_prefetchable                   ("false"),
		.vendor_id                           (4466),
		.device_id                           (57345),
		.revision_id                         (1),
		.class_code                          (0),
		.subsystem_vendor_id                 (4466),
		.subsystem_device_id                 (4),
		.port_link_number                    (1),
		.msi_function_count                  (0),
		.enable_msi_64bit_addressing         ("true"),
		.enable_function_msix_support        ("false"),
		.eie_before_nfts_count               (4),
		.enable_completion_timeout_disable   ("false"),
		.completion_timeout                  ("NONE"),
		.enable_adapter_half_rate_mode       ("false"),
		.msix_pba_bir                        (0),
		.msix_pba_offset                     (0),
		.msix_table_bir                      (0),
		.msix_table_offset                   (0),
		.msix_table_size                     (0),
		.use_crc_forwarding                  ("false"),
		.surprise_down_error_support         ("false"),
		.dll_active_report_support           ("false"),
		.bar_io_window_size                  ("32BIT"),
		.bar_prefetchable                    (32),
		.hot_plug_support                    (7'b0000000),
		.no_command_completed                ("true"),
		.slot_power_limit                    (0),
		.slot_power_scale                    (0),
		.slot_number                         (0),
		.enable_slot_register                ("false"),
		.advanced_errors                     ("false"),
		.enable_ecrc_check                   ("false"),
		.enable_ecrc_gen                     ("false"),
		.max_payload_size                    (0),
		.retry_buffer_last_active_address    (255),
		.credit_buffer_allocation_aux        ("ABSOLUTE"),
		.vc0_rx_flow_ctrl_posted_header      (28),
		.vc0_rx_flow_ctrl_posted_data        (198),
		.vc0_rx_flow_ctrl_nonposted_header   (30),
		.vc0_rx_flow_ctrl_nonposted_data     (0),
		.vc0_rx_flow_ctrl_compl_header       (48),
		.vc0_rx_flow_ctrl_compl_data         (256),
		.RX_BUF                              (9),
		.RH_NUM                              (7),
		.G_TAG_NUM0                          (32),
		.endpoint_l0_latency                 (0),
		.endpoint_l1_latency                 (0),
		.enable_l1_aspm                      ("false"),
		.l01_entry_latency                   (31),
		.diffclock_nfts_count                (255),
		.sameclock_nfts_count                (255),
		.l1_exit_latency_sameclock           (7),
		.l1_exit_latency_diffclock           (7),
		.l0_exit_latency_sameclock           (7),
		.l0_exit_latency_diffclock           (7),
		.gen2_diffclock_nfts_count           (255),
		.gen2_sameclock_nfts_count           (255),
		.CG_COMMON_CLOCK_MODE                (1),
		.CB_PCIE_MODE                        (0),
		.AST_LITE                            (0),
		.CB_PCIE_RX_LITE                     (0),
		.CG_RXM_IRQ_NUM                      (16),
		.CG_AVALON_S_ADDR_WIDTH              (20),
		.bypass_tl                           ("false"),
		.CG_IMPL_CRA_AV_SLAVE_PORT           (1),
		.CG_NO_CPL_REORDERING                (0),
		.CG_ENABLE_A2P_INTERRUPT             (0),
		.p_user_msi_enable                   (0),
		.CG_IRQ_BIT_ENA                      (65535),
		.CB_A2P_ADDR_MAP_IS_FIXED            (1),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES         (1),
		.CB_A2P_ADDR_MAP_PASS_THRU_BITS      (31),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_LOW  (32'b00000000000000000000000000000000),
		.RXM_DATA_WIDTH                      (64),
		.RXM_BEN_WIDTH                       (8),
		.TL_SELECTION                        (1),
		.pcie_mode                           ("SHARED_MODE"),
		.single_rx_detect                    (1),
		.enable_coreclk_out_half_rate        ("false"),
		.low_priority_vc                     (0),
		.link_width                          (1),
		.cyclone4                            (1)
	) pcie_ip (
		.pcie_core_clk_clk                  (pcie_ip_pcie_core_clk_clk),                   //      pcie_core_clk.clk
		.pcie_core_reset_reset_n            (pcie_ip_pcie_core_reset_reset),               //    pcie_core_reset.reset_n
		.cal_blk_clk_clk                    (altpll_qsys_c3_clk),                          //        cal_blk_clk.clk
		.txs_address                        (mm_interconnect_1_pcie_ip_txs_address),       //                txs.address
		.txs_chipselect                     (mm_interconnect_1_pcie_ip_txs_chipselect),    //                   .chipselect
		.txs_byteenable                     (mm_interconnect_1_pcie_ip_txs_byteenable),    //                   .byteenable
		.txs_readdata                       (mm_interconnect_1_pcie_ip_txs_readdata),      //                   .readdata
		.txs_writedata                      (mm_interconnect_1_pcie_ip_txs_writedata),     //                   .writedata
		.txs_read                           (mm_interconnect_1_pcie_ip_txs_read),          //                   .read
		.txs_write                          (mm_interconnect_1_pcie_ip_txs_write),         //                   .write
		.txs_burstcount                     (mm_interconnect_1_pcie_ip_txs_burstcount),    //                   .burstcount
		.txs_readdatavalid                  (mm_interconnect_1_pcie_ip_txs_readdatavalid), //                   .readdatavalid
		.txs_waitrequest                    (mm_interconnect_1_pcie_ip_txs_waitrequest),   //                   .waitrequest
		.refclk_export                      (pcie_ip_refclk_export),                       //             refclk.export
		.test_in_test_in                    (pcie_ip_test_in_test_in),                     //            test_in.test_in
		.pcie_rstn_export                   (pcie_ip_pcie_rstn_export),                    //          pcie_rstn.export
		.clocks_sim_clk250_export           (pcie_ip_clocks_sim_clk250_export),            //         clocks_sim.clk250_export
		.clocks_sim_clk500_export           (pcie_ip_clocks_sim_clk500_export),            //                   .clk500_export
		.clocks_sim_clk125_export           (pcie_ip_clocks_sim_clk125_export),            //                   .clk125_export
		.reconfig_busy_busy_altgxb_reconfig (pcie_ip_reconfig_busy_busy_altgxb_reconfig),  //      reconfig_busy.busy_altgxb_reconfig
		.pipe_ext_pipe_mode                 (pcie_ip_pipe_ext_pipe_mode),                  //           pipe_ext.pipe_mode
		.pipe_ext_phystatus_ext             (pcie_ip_pipe_ext_phystatus_ext),              //                   .phystatus_ext
		.pipe_ext_rate_ext                  (pcie_ip_pipe_ext_rate_ext),                   //                   .rate_ext
		.pipe_ext_powerdown_ext             (pcie_ip_pipe_ext_powerdown_ext),              //                   .powerdown_ext
		.pipe_ext_txdetectrx_ext            (pcie_ip_pipe_ext_txdetectrx_ext),             //                   .txdetectrx_ext
		.pipe_ext_rxelecidle0_ext           (pcie_ip_pipe_ext_rxelecidle0_ext),            //                   .rxelecidle0_ext
		.pipe_ext_rxdata0_ext               (pcie_ip_pipe_ext_rxdata0_ext),                //                   .rxdata0_ext
		.pipe_ext_rxstatus0_ext             (pcie_ip_pipe_ext_rxstatus0_ext),              //                   .rxstatus0_ext
		.pipe_ext_rxvalid0_ext              (pcie_ip_pipe_ext_rxvalid0_ext),               //                   .rxvalid0_ext
		.pipe_ext_rxdatak0_ext              (pcie_ip_pipe_ext_rxdatak0_ext),               //                   .rxdatak0_ext
		.pipe_ext_txdata0_ext               (pcie_ip_pipe_ext_txdata0_ext),                //                   .txdata0_ext
		.pipe_ext_txdatak0_ext              (pcie_ip_pipe_ext_txdatak0_ext),               //                   .txdatak0_ext
		.pipe_ext_rxpolarity0_ext           (pcie_ip_pipe_ext_rxpolarity0_ext),            //                   .rxpolarity0_ext
		.pipe_ext_txcompl0_ext              (pcie_ip_pipe_ext_txcompl0_ext),               //                   .txcompl0_ext
		.pipe_ext_txelecidle0_ext           (pcie_ip_pipe_ext_txelecidle0_ext),            //                   .txelecidle0_ext
		.powerdown_pll_powerdown            (pcie_ip_powerdown_pll_powerdown),             //          powerdown.pll_powerdown
		.powerdown_gxb_powerdown            (pcie_ip_powerdown_gxb_powerdown),             //                   .gxb_powerdown
		.bar1_0_address                     (pcie_ip_bar1_0_address),                      //             bar1_0.address
		.bar1_0_read                        (pcie_ip_bar1_0_read),                         //                   .read
		.bar1_0_waitrequest                 (pcie_ip_bar1_0_waitrequest),                  //                   .waitrequest
		.bar1_0_write                       (pcie_ip_bar1_0_write),                        //                   .write
		.bar1_0_readdatavalid               (pcie_ip_bar1_0_readdatavalid),                //                   .readdatavalid
		.bar1_0_readdata                    (pcie_ip_bar1_0_readdata),                     //                   .readdata
		.bar1_0_writedata                   (pcie_ip_bar1_0_writedata),                    //                   .writedata
		.bar1_0_burstcount                  (pcie_ip_bar1_0_burstcount),                   //                   .burstcount
		.bar1_0_byteenable                  (pcie_ip_bar1_0_byteenable),                   //                   .byteenable
		.bar2_address                       (pcie_ip_bar2_address),                        //               bar2.address
		.bar2_read                          (pcie_ip_bar2_read),                           //                   .read
		.bar2_waitrequest                   (pcie_ip_bar2_waitrequest),                    //                   .waitrequest
		.bar2_write                         (pcie_ip_bar2_write),                          //                   .write
		.bar2_readdatavalid                 (pcie_ip_bar2_readdatavalid),                  //                   .readdatavalid
		.bar2_readdata                      (pcie_ip_bar2_readdata),                       //                   .readdata
		.bar2_writedata                     (pcie_ip_bar2_writedata),                      //                   .writedata
		.bar2_burstcount                    (pcie_ip_bar2_burstcount),                     //                   .burstcount
		.bar2_byteenable                    (pcie_ip_bar2_byteenable),                     //                   .byteenable
		.cra_chipselect                     (mm_interconnect_0_pcie_ip_cra_chipselect),    //                cra.chipselect
		.cra_address                        (mm_interconnect_0_pcie_ip_cra_address),       //                   .address
		.cra_byteenable                     (mm_interconnect_0_pcie_ip_cra_byteenable),    //                   .byteenable
		.cra_read                           (mm_interconnect_0_pcie_ip_cra_read),          //                   .read
		.cra_readdata                       (mm_interconnect_0_pcie_ip_cra_readdata),      //                   .readdata
		.cra_write                          (mm_interconnect_0_pcie_ip_cra_write),         //                   .write
		.cra_writedata                      (mm_interconnect_0_pcie_ip_cra_writedata),     //                   .writedata
		.cra_waitrequest                    (mm_interconnect_0_pcie_ip_cra_waitrequest),   //                   .waitrequest
		.cra_irq_irq                        (),                                            //            cra_irq.irq
		.rxm_irq_irq                        (pcie_ip_rxm_irq_irq),                         //            rxm_irq.irq
		.rx_in_rx_datain_0                  (pcie_ip_rx_in_rx_datain_0),                   //              rx_in.rx_datain_0
		.tx_out_tx_dataout_0                (pcie_ip_tx_out_tx_dataout_0),                 //             tx_out.tx_dataout_0
		.reconfig_togxb_data                (pcie_ip_reconfig_togxb_data),                 //     reconfig_togxb.data
		.reconfig_gxbclk_clk                (altpll_qsys_c3_clk),                          //    reconfig_gxbclk.clk
		.reconfig_fromgxb_0_data            (pcie_ip_reconfig_fromgxb_0_data),             // reconfig_fromgxb_0.data
		.fixedclk_clk                       (pcie_ip_pcie_core_clk_clk)                    //           fixedclk.clk
	);

	ahb_master_slave_with_pcie_sgdma sgdma (
		.clk                           (pcie_ip_pcie_core_clk_clk),              //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),        //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),               //          csr_irq.irq
		.m_read_readdata               (sgdma_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_m_read_read),                      //                 .read
		.m_read_burstcount             (sgdma_m_read_burstcount),                //                 .burstcount
		.m_write_waitrequest           (sgdma_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_m_write_byteenable),               //                 .byteenable
		.m_write_burstcount            (sgdma_m_write_burstcount)                //                 .burstcount
	);

	ahb_master_slave_with_pcie_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	ahb_master_slave_with_pcie_altpll_qsys altpll_qsys (
		.clk       (clk_clk),                            //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                                   //             pll_slave.read
		.write     (),                                   //                      .write
		.address   (),                                   //                      .address
		.readdata  (),                                   //                      .readdata
		.writedata (),                                   //                      .writedata
		.c0        (),                                   //                    c0.clk
		.c1        (altpll_sdram_clk),                   //                    c1.clk
		.c2        (),                                   //                    c2.clk
		.c3        (altpll_qsys_c3_clk),                 //                    c3.clk
		.areset    (),                                   //        areset_conduit.export
		.locked    (),                                   //        locked_conduit.export
		.phasedone ()                                    //     phasedone_conduit.export
	);

	avalon_ahb_bridge #(
		.AVALON_ADDRESSWIDTH (5),
		.ADDRESSWIDTH        (32),
		.DATAWIDTH           (32)
	) avalon2ahb_bridge_0 (
		.clk           (clk_clk),                                                          //        clock.clk
		.reset_n       (~rst_controller_002_reset_out_reset),                              //        reset.reset_n
		.read          (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_read),          // avalon_slave.read
		.address       (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_address),       //             .address
		.write         (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_write),         //             .write
		.writedata     (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_writedata),     //             .writedata
		.waitrequest   (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_waitrequest),   //             .waitrequest
		.readdatavalid (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_readdatavalid), //             .readdatavalid
		.readdata      (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_readdata),      //             .readdata
		.HRDATA        (avalon2ahb_bridge_0_ahb_master_hrdata),                            //   ahb_master.hrdata
		.HREADY        (avalon2ahb_bridge_0_ahb_master_hready),                            //             .hready
		.HRESP         (avalon2ahb_bridge_0_ahb_master_hresp),                             //             .hresp
		.HBURST        (avalon2ahb_bridge_0_ahb_master_hburst),                            //             .hburst
		.HSIZE         (avalon2ahb_bridge_0_ahb_master_hsize),                             //             .hsize
		.HTRANS        (avalon2ahb_bridge_0_ahb_master_htrans),                            //             .htrans
		.HSEL          (avalon2ahb_bridge_0_ahb_master_hsel),                              //             .hsel
		.HPROT         (avalon2ahb_bridge_0_ahb_master_hprot),                             //             .hprot
		.HADDR         (avalon2ahb_bridge_0_ahb_master_haddr),                             //             .haddr
		.HWDATA        (avalon2ahb_bridge_0_ahb_master_hwdata),                            //             .hwdata
		.HWRITE        (avalon2ahb_bridge_0_ahb_master_hwrite),                            //             .hwrite
		.HREADYIN      (avalon2ahb_bridge_0_ahb_master_hreadyin)                           //             .hreadyin
	);

	top_level ahb_master_slave_2_0 (
		.add_data_sel    (ahb_master_slave_2_0_conduit_end_add_data_sel), // conduit_end.add_data_sel
		.rdwr_address    (ahb_master_slave_2_0_conduit_end_rdwr_address), //            .rdwr_address
		.display_data    (ahb_master_slave_2_0_conduit_end_display_data), //            .display_data
		.HRESETn         (~rst_controller_002_reset_out_reset),           //  reset_sink.reset_n
		.HCLK            (clk_clk),                                       //  clock_sink.clk
		.slave_HADDR     (avalon2ahb_bridge_0_ahb_master_haddr),          //   ahb_slave.haddr
		.slave_HBURST    (avalon2ahb_bridge_0_ahb_master_hburst),         //            .hburst
		.slave_HPROT     (avalon2ahb_bridge_0_ahb_master_hprot),          //            .hprot
		.slave_HSIZE     (avalon2ahb_bridge_0_ahb_master_hsize),          //            .hsize
		.slave_HTRANS    (avalon2ahb_bridge_0_ahb_master_htrans),         //            .htrans
		.slave_HWDATA    (avalon2ahb_bridge_0_ahb_master_hwdata),         //            .hwdata
		.slave_HWRITE    (avalon2ahb_bridge_0_ahb_master_hwrite),         //            .hwrite
		.slave_HRDATA    (avalon2ahb_bridge_0_ahb_master_hrdata),         //            .hrdata
		.slave_HREADYOUT (avalon2ahb_bridge_0_ahb_master_hready),         //            .hready
		.slave_HRESP     (avalon2ahb_bridge_0_ahb_master_hresp),          //            .hresp
		.slave_HSEL      (avalon2ahb_bridge_0_ahb_master_hsel),           //            .hsel
		.slave_HREADY    (avalon2ahb_bridge_0_ahb_master_hreadyin),       //            .hreadyin
		.master_HADDR    (ahb_master_slave_2_0_ahb_master_haddr),         //  ahb_master.haddr
		.master_HBURST   (ahb_master_slave_2_0_ahb_master_hburst),        //            .hburst
		.master_HPROT    (ahb_master_slave_2_0_ahb_master_hprot),         //            .hprot
		.master_HSIZE    (ahb_master_slave_2_0_ahb_master_hsize),         //            .hsize
		.master_HTRANS   (ahb_master_slave_2_0_ahb_master_htrans),        //            .htrans
		.master_HWDATA   (ahb_master_slave_2_0_ahb_master_hwdata),        //            .hwdata
		.master_HWRITE   (ahb_master_slave_2_0_ahb_master_hwrite),        //            .hwrite
		.master_HRDATA   (ahb_master_slave_2_0_ahb_master_hrdata),        //            .hrdata
		.master_HREADY   (ahb_master_slave_2_0_ahb_master_hready),        //            .hready
		.master_HRESP    (ahb_master_slave_2_0_ahb_master_hresp),         //            .hresp
		.master_HREADYIN (ahb_master_slave_2_0_ahb_master_hreadyin),      //            .hreadyin
		.master_HSEL     (ahb_master_slave_2_0_ahb_master_hsel)           //            .hsel
	);

	ahb_avalon_bridge_with_burst #(
		.ADDRESSWIDTH  (32),
		.DATAWIDTH     (32),
		.FIFODEPTH     (32),
		.FIFODEPTH_LOG (5),
		.MAXBURSTCOUNT (8)
	) ahb2avalon_burst_bridge_0 (
		.clk           (clk_clk),                                               //         clock.clk
		.reset_n       (~rst_controller_002_reset_out_reset),                   //         reset.reset_n
		.address       (ahb2avalon_burst_bridge_0_avalon_master_address),       // avalon_master.address
		.write         (ahb2avalon_burst_bridge_0_avalon_master_write),         //              .write
		.read          (ahb2avalon_burst_bridge_0_avalon_master_read),          //              .read
		.byteenable    (ahb2avalon_burst_bridge_0_avalon_master_byteenable),    //              .byteenable
		.writedata     (ahb2avalon_burst_bridge_0_avalon_master_writedata),     //              .writedata
		.waitrequest   (ahb2avalon_burst_bridge_0_avalon_master_waitrequest),   //              .waitrequest
		.readdatavalid (ahb2avalon_burst_bridge_0_avalon_master_readdatavalid), //              .readdatavalid
		.readdata      (ahb2avalon_burst_bridge_0_avalon_master_readdata),      //              .readdata
		.burstcount    (ahb2avalon_burst_bridge_0_avalon_master_burstcount),    //              .burstcount
		.HRDATA        (ahb_master_slave_2_0_ahb_master_hrdata),                //     ahb_slave.hrdata
		.HREADY        (ahb_master_slave_2_0_ahb_master_hreadyin),              //              .hreadyin
		.HRESP         (ahb_master_slave_2_0_ahb_master_hresp),                 //              .hresp
		.HBURST        (ahb_master_slave_2_0_ahb_master_hburst),                //              .hburst
		.HSIZE         (ahb_master_slave_2_0_ahb_master_hsize),                 //              .hsize
		.HTRANS        (ahb_master_slave_2_0_ahb_master_htrans),                //              .htrans
		.HPROT         (ahb_master_slave_2_0_ahb_master_hprot),                 //              .hprot
		.HADDR         (ahb_master_slave_2_0_ahb_master_haddr),                 //              .haddr
		.HWDATA        (ahb_master_slave_2_0_ahb_master_hwdata),                //              .hwdata
		.HWRITE        (ahb_master_slave_2_0_ahb_master_hwrite),                //              .hwrite
		.HREADYOUT     (ahb_master_slave_2_0_ahb_master_hready),                //              .hready
		.HSEL          (ahb_master_slave_2_0_ahb_master_hsel)                   //              .hsel
	);

	ahb_master_slave_with_pcie_mm_interconnect_0 mm_interconnect_0 (
		.pcie_ip_pcie_core_clk_clk                                 (pcie_ip_pcie_core_clk_clk),                 //                               pcie_ip_pcie_core_clk.clk
		.pcie_ip_bar2_translator_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),        // pcie_ip_bar2_translator_reset_reset_bridge_in_reset.reset
		.sgdma_reset_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),            //                   sgdma_reset_reset_bridge_in_reset.reset
		.pcie_ip_bar2_address                                      (pcie_ip_bar2_address),                      //                                        pcie_ip_bar2.address
		.pcie_ip_bar2_waitrequest                                  (pcie_ip_bar2_waitrequest),                  //                                                    .waitrequest
		.pcie_ip_bar2_burstcount                                   (pcie_ip_bar2_burstcount),                   //                                                    .burstcount
		.pcie_ip_bar2_byteenable                                   (pcie_ip_bar2_byteenable),                   //                                                    .byteenable
		.pcie_ip_bar2_read                                         (pcie_ip_bar2_read),                         //                                                    .read
		.pcie_ip_bar2_readdata                                     (pcie_ip_bar2_readdata),                     //                                                    .readdata
		.pcie_ip_bar2_readdatavalid                                (pcie_ip_bar2_readdatavalid),                //                                                    .readdatavalid
		.pcie_ip_bar2_write                                        (pcie_ip_bar2_write),                        //                                                    .write
		.pcie_ip_bar2_writedata                                    (pcie_ip_bar2_writedata),                    //                                                    .writedata
		.pcie_ip_cra_address                                       (mm_interconnect_0_pcie_ip_cra_address),     //                                         pcie_ip_cra.address
		.pcie_ip_cra_write                                         (mm_interconnect_0_pcie_ip_cra_write),       //                                                    .write
		.pcie_ip_cra_read                                          (mm_interconnect_0_pcie_ip_cra_read),        //                                                    .read
		.pcie_ip_cra_readdata                                      (mm_interconnect_0_pcie_ip_cra_readdata),    //                                                    .readdata
		.pcie_ip_cra_writedata                                     (mm_interconnect_0_pcie_ip_cra_writedata),   //                                                    .writedata
		.pcie_ip_cra_byteenable                                    (mm_interconnect_0_pcie_ip_cra_byteenable),  //                                                    .byteenable
		.pcie_ip_cra_waitrequest                                   (mm_interconnect_0_pcie_ip_cra_waitrequest), //                                                    .waitrequest
		.pcie_ip_cra_chipselect                                    (mm_interconnect_0_pcie_ip_cra_chipselect),  //                                                    .chipselect
		.sgdma_csr_address                                         (mm_interconnect_0_sgdma_csr_address),       //                                           sgdma_csr.address
		.sgdma_csr_write                                           (mm_interconnect_0_sgdma_csr_write),         //                                                    .write
		.sgdma_csr_read                                            (mm_interconnect_0_sgdma_csr_read),          //                                                    .read
		.sgdma_csr_readdata                                        (mm_interconnect_0_sgdma_csr_readdata),      //                                                    .readdata
		.sgdma_csr_writedata                                       (mm_interconnect_0_sgdma_csr_writedata),     //                                                    .writedata
		.sgdma_csr_chipselect                                      (mm_interconnect_0_sgdma_csr_chipselect)     //                                                    .chipselect
	);

	ahb_master_slave_with_pcie_mm_interconnect_1 mm_interconnect_1 (
		.clk_50_clk_clk                                              (clk_clk),                                               //                                            clk_50_clk.clk
		.pcie_ip_pcie_core_clk_clk                                   (pcie_ip_pcie_core_clk_clk),                             //                                 pcie_ip_pcie_core_clk.clk
		.ahb2avalon_burst_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                    // ahb2avalon_burst_bridge_0_reset_reset_bridge_in_reset.reset
		.pcie_ip_txs_translator_reset_reset_bridge_in_reset_reset    (rst_controller_003_reset_out_reset),                    //    pcie_ip_txs_translator_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset                     (rst_controller_001_reset_out_reset),                    //                     sdram_reset_reset_bridge_in_reset.reset
		.sgdma_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                        //                     sgdma_reset_reset_bridge_in_reset.reset
		.ahb2avalon_burst_bridge_0_avalon_master_address             (ahb2avalon_burst_bridge_0_avalon_master_address),       //               ahb2avalon_burst_bridge_0_avalon_master.address
		.ahb2avalon_burst_bridge_0_avalon_master_waitrequest         (ahb2avalon_burst_bridge_0_avalon_master_waitrequest),   //                                                      .waitrequest
		.ahb2avalon_burst_bridge_0_avalon_master_burstcount          (ahb2avalon_burst_bridge_0_avalon_master_burstcount),    //                                                      .burstcount
		.ahb2avalon_burst_bridge_0_avalon_master_byteenable          (ahb2avalon_burst_bridge_0_avalon_master_byteenable),    //                                                      .byteenable
		.ahb2avalon_burst_bridge_0_avalon_master_read                (ahb2avalon_burst_bridge_0_avalon_master_read),          //                                                      .read
		.ahb2avalon_burst_bridge_0_avalon_master_readdata            (ahb2avalon_burst_bridge_0_avalon_master_readdata),      //                                                      .readdata
		.ahb2avalon_burst_bridge_0_avalon_master_readdatavalid       (ahb2avalon_burst_bridge_0_avalon_master_readdatavalid), //                                                      .readdatavalid
		.ahb2avalon_burst_bridge_0_avalon_master_write               (ahb2avalon_burst_bridge_0_avalon_master_write),         //                                                      .write
		.ahb2avalon_burst_bridge_0_avalon_master_writedata           (ahb2avalon_burst_bridge_0_avalon_master_writedata),     //                                                      .writedata
		.sgdma_descriptor_read_address                               (sgdma_descriptor_read_address),                         //                                 sgdma_descriptor_read.address
		.sgdma_descriptor_read_waitrequest                           (sgdma_descriptor_read_waitrequest),                     //                                                      .waitrequest
		.sgdma_descriptor_read_read                                  (sgdma_descriptor_read_read),                            //                                                      .read
		.sgdma_descriptor_read_readdata                              (sgdma_descriptor_read_readdata),                        //                                                      .readdata
		.sgdma_descriptor_read_readdatavalid                         (sgdma_descriptor_read_readdatavalid),                   //                                                      .readdatavalid
		.sgdma_descriptor_write_address                              (sgdma_descriptor_write_address),                        //                                sgdma_descriptor_write.address
		.sgdma_descriptor_write_waitrequest                          (sgdma_descriptor_write_waitrequest),                    //                                                      .waitrequest
		.sgdma_descriptor_write_write                                (sgdma_descriptor_write_write),                          //                                                      .write
		.sgdma_descriptor_write_writedata                            (sgdma_descriptor_write_writedata),                      //                                                      .writedata
		.sgdma_m_read_address                                        (sgdma_m_read_address),                                  //                                          sgdma_m_read.address
		.sgdma_m_read_waitrequest                                    (sgdma_m_read_waitrequest),                              //                                                      .waitrequest
		.sgdma_m_read_burstcount                                     (sgdma_m_read_burstcount),                               //                                                      .burstcount
		.sgdma_m_read_read                                           (sgdma_m_read_read),                                     //                                                      .read
		.sgdma_m_read_readdata                                       (sgdma_m_read_readdata),                                 //                                                      .readdata
		.sgdma_m_read_readdatavalid                                  (sgdma_m_read_readdatavalid),                            //                                                      .readdatavalid
		.sgdma_m_write_address                                       (sgdma_m_write_address),                                 //                                         sgdma_m_write.address
		.sgdma_m_write_waitrequest                                   (sgdma_m_write_waitrequest),                             //                                                      .waitrequest
		.sgdma_m_write_burstcount                                    (sgdma_m_write_burstcount),                              //                                                      .burstcount
		.sgdma_m_write_byteenable                                    (sgdma_m_write_byteenable),                              //                                                      .byteenable
		.sgdma_m_write_write                                         (sgdma_m_write_write),                                   //                                                      .write
		.sgdma_m_write_writedata                                     (sgdma_m_write_writedata),                               //                                                      .writedata
		.pcie_ip_txs_address                                         (mm_interconnect_1_pcie_ip_txs_address),                 //                                           pcie_ip_txs.address
		.pcie_ip_txs_write                                           (mm_interconnect_1_pcie_ip_txs_write),                   //                                                      .write
		.pcie_ip_txs_read                                            (mm_interconnect_1_pcie_ip_txs_read),                    //                                                      .read
		.pcie_ip_txs_readdata                                        (mm_interconnect_1_pcie_ip_txs_readdata),                //                                                      .readdata
		.pcie_ip_txs_writedata                                       (mm_interconnect_1_pcie_ip_txs_writedata),               //                                                      .writedata
		.pcie_ip_txs_burstcount                                      (mm_interconnect_1_pcie_ip_txs_burstcount),              //                                                      .burstcount
		.pcie_ip_txs_byteenable                                      (mm_interconnect_1_pcie_ip_txs_byteenable),              //                                                      .byteenable
		.pcie_ip_txs_readdatavalid                                   (mm_interconnect_1_pcie_ip_txs_readdatavalid),           //                                                      .readdatavalid
		.pcie_ip_txs_waitrequest                                     (mm_interconnect_1_pcie_ip_txs_waitrequest),             //                                                      .waitrequest
		.pcie_ip_txs_chipselect                                      (mm_interconnect_1_pcie_ip_txs_chipselect),              //                                                      .chipselect
		.sdram_s1_address                                            (mm_interconnect_1_sdram_s1_address),                    //                                              sdram_s1.address
		.sdram_s1_write                                              (mm_interconnect_1_sdram_s1_write),                      //                                                      .write
		.sdram_s1_read                                               (mm_interconnect_1_sdram_s1_read),                       //                                                      .read
		.sdram_s1_readdata                                           (mm_interconnect_1_sdram_s1_readdata),                   //                                                      .readdata
		.sdram_s1_writedata                                          (mm_interconnect_1_sdram_s1_writedata),                  //                                                      .writedata
		.sdram_s1_byteenable                                         (mm_interconnect_1_sdram_s1_byteenable),                 //                                                      .byteenable
		.sdram_s1_readdatavalid                                      (mm_interconnect_1_sdram_s1_readdatavalid),              //                                                      .readdatavalid
		.sdram_s1_waitrequest                                        (mm_interconnect_1_sdram_s1_waitrequest),                //                                                      .waitrequest
		.sdram_s1_chipselect                                         (mm_interconnect_1_sdram_s1_chipselect)                  //                                                      .chipselect
	);

	ahb_master_slave_with_pcie_mm_interconnect_2 mm_interconnect_2 (
		.clk_50_clk_clk                                              (clk_clk),                                                          //                                            clk_50_clk.clk
		.pcie_ip_pcie_core_clk_clk                                   (pcie_ip_pcie_core_clk_clk),                                        //                                 pcie_ip_pcie_core_clk.clk
		.avalon2ahb_bridge_0_reset_reset_bridge_in_reset_reset       (rst_controller_002_reset_out_reset),                               //       avalon2ahb_bridge_0_reset_reset_bridge_in_reset.reset
		.pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                               // pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset.reset
		.pcie_ip_bar1_0_address                                      (pcie_ip_bar1_0_address),                                           //                                        pcie_ip_bar1_0.address
		.pcie_ip_bar1_0_waitrequest                                  (pcie_ip_bar1_0_waitrequest),                                       //                                                      .waitrequest
		.pcie_ip_bar1_0_burstcount                                   (pcie_ip_bar1_0_burstcount),                                        //                                                      .burstcount
		.pcie_ip_bar1_0_byteenable                                   (pcie_ip_bar1_0_byteenable),                                        //                                                      .byteenable
		.pcie_ip_bar1_0_read                                         (pcie_ip_bar1_0_read),                                              //                                                      .read
		.pcie_ip_bar1_0_readdata                                     (pcie_ip_bar1_0_readdata),                                          //                                                      .readdata
		.pcie_ip_bar1_0_readdatavalid                                (pcie_ip_bar1_0_readdatavalid),                                     //                                                      .readdatavalid
		.pcie_ip_bar1_0_write                                        (pcie_ip_bar1_0_write),                                             //                                                      .write
		.pcie_ip_bar1_0_writedata                                    (pcie_ip_bar1_0_writedata),                                         //                                                      .writedata
		.avalon2ahb_bridge_0_avalon_slave_address                    (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_address),       //                      avalon2ahb_bridge_0_avalon_slave.address
		.avalon2ahb_bridge_0_avalon_slave_write                      (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_write),         //                                                      .write
		.avalon2ahb_bridge_0_avalon_slave_read                       (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_read),          //                                                      .read
		.avalon2ahb_bridge_0_avalon_slave_readdata                   (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_readdata),      //                                                      .readdata
		.avalon2ahb_bridge_0_avalon_slave_writedata                  (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_writedata),     //                                                      .writedata
		.avalon2ahb_bridge_0_avalon_slave_readdatavalid              (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_readdatavalid), //                                                      .readdatavalid
		.avalon2ahb_bridge_0_avalon_slave_waitrequest                (mm_interconnect_2_avalon2ahb_bridge_0_avalon_slave_waitrequest)    //                                                      .waitrequest
	);

	ahb_master_slave_with_pcie_irq_mapper irq_mapper (
		.clk           (pcie_ip_pcie_core_clk_clk),          //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (pcie_ip_rxm_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.reset_in1      (~pcie_ip_pcie_core_reset_reset), // reset_in1.reset
		.clk            (pcie_ip_pcie_core_clk_clk),      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~pcie_ip_pcie_core_reset_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~pcie_ip_pcie_core_reset_reset),     // reset_in0.reset
		.clk            (pcie_ip_pcie_core_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
