library verilog;
use verilog.vl_types.all;
entity verbosity_pkg is
end verbosity_pkg;
