library verilog;
use verilog.vl_types.all;
entity ama_multiplier_function is
    generic(
        width_data_in_a : integer := 1;
        width_data_in_b : integer := 1;
        width_data_out  : integer := 1;
        number_of_multipliers: integer := 1;
        multiplier_input_representation_a: string  := "UNSIGNED";
        multiplier_input_representation_b: string  := "UNSIGNED";
        multiplier_register0: string  := "UNREGISTERED";
        multiplier_register1: string  := "UNREGISTERED";
        multiplier_register2: string  := "UNREGISTERED";
        multiplier_register3: string  := "UNREGISTERED";
        multiplier_aclr0: string  := "NONE";
        multiplier_aclr1: string  := "NONE";
        multiplier_aclr2: string  := "NONE";
        multiplier_aclr3: string  := "NONE";
        width_data_in_a_msb: vl_notype;
        width_data_in_b_msb: vl_notype;
        width_data_out_msb: vl_notype;
        width_mult_input_a: vl_notype;
        width_mult_input_a_msb: vl_notype;
        width_mult_input_b: vl_notype;
        width_mult_input_b_msb: vl_notype;
        width_mult_output: vl_notype
    );
    port(
        clock           : in     vl_logic_vector(3 downto 0);
        aclr            : in     vl_logic_vector(3 downto 0);
        ena             : in     vl_logic_vector(3 downto 0);
        data_in_a0      : in     vl_logic_vector;
        data_in_a1      : in     vl_logic_vector;
        data_in_a2      : in     vl_logic_vector;
        data_in_a3      : in     vl_logic_vector;
        data_in_b0      : in     vl_logic_vector;
        data_in_b1      : in     vl_logic_vector;
        data_in_b2      : in     vl_logic_vector;
        data_in_b3      : in     vl_logic_vector;
        data_out_0      : out    vl_logic_vector;
        data_out_1      : out    vl_logic_vector;
        data_out_2      : out    vl_logic_vector;
        data_out_3      : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of width_data_in_a : constant is 1;
    attribute mti_svvh_generic_type of width_data_in_b : constant is 1;
    attribute mti_svvh_generic_type of width_data_out : constant is 1;
    attribute mti_svvh_generic_type of number_of_multipliers : constant is 1;
    attribute mti_svvh_generic_type of multiplier_input_representation_a : constant is 1;
    attribute mti_svvh_generic_type of multiplier_input_representation_b : constant is 1;
    attribute mti_svvh_generic_type of multiplier_register0 : constant is 1;
    attribute mti_svvh_generic_type of multiplier_register1 : constant is 1;
    attribute mti_svvh_generic_type of multiplier_register2 : constant is 1;
    attribute mti_svvh_generic_type of multiplier_register3 : constant is 1;
    attribute mti_svvh_generic_type of multiplier_aclr0 : constant is 1;
    attribute mti_svvh_generic_type of multiplier_aclr1 : constant is 1;
    attribute mti_svvh_generic_type of multiplier_aclr2 : constant is 1;
    attribute mti_svvh_generic_type of multiplier_aclr3 : constant is 1;
    attribute mti_svvh_generic_type of width_data_in_a_msb : constant is 3;
    attribute mti_svvh_generic_type of width_data_in_b_msb : constant is 3;
    attribute mti_svvh_generic_type of width_data_out_msb : constant is 3;
    attribute mti_svvh_generic_type of width_mult_input_a : constant is 3;
    attribute mti_svvh_generic_type of width_mult_input_a_msb : constant is 3;
    attribute mti_svvh_generic_type of width_mult_input_b : constant is 3;
    attribute mti_svvh_generic_type of width_mult_input_b_msb : constant is 3;
    attribute mti_svvh_generic_type of width_mult_output : constant is 3;
end ama_multiplier_function;
