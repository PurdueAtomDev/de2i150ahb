library verilog;
use verilog.vl_types.all;
entity avalon_mm_pkg is
end avalon_mm_pkg;
